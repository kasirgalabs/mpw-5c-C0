magic
tech sky130A
magscale 1 2
timestamp 1647257906
<< obsli1 >>
rect 1104 2159 258888 257329
<< obsm1 >>
rect 566 1980 258888 257360
<< metal2 >>
rect 1674 0 1730 800
rect 5078 0 5134 800
rect 8574 0 8630 800
rect 12070 0 12126 800
rect 15474 0 15530 800
rect 18970 0 19026 800
rect 22466 0 22522 800
rect 25870 0 25926 800
rect 29366 0 29422 800
rect 32862 0 32918 800
rect 36266 0 36322 800
rect 39762 0 39818 800
rect 43258 0 43314 800
rect 46662 0 46718 800
rect 50158 0 50214 800
rect 53654 0 53710 800
rect 57058 0 57114 800
rect 60554 0 60610 800
rect 64050 0 64106 800
rect 67454 0 67510 800
rect 70950 0 71006 800
rect 74446 0 74502 800
rect 77850 0 77906 800
rect 81346 0 81402 800
rect 84842 0 84898 800
rect 88338 0 88394 800
rect 91742 0 91798 800
rect 95238 0 95294 800
rect 98734 0 98790 800
rect 102138 0 102194 800
rect 105634 0 105690 800
rect 109130 0 109186 800
rect 112534 0 112590 800
rect 116030 0 116086 800
rect 119526 0 119582 800
rect 122930 0 122986 800
rect 126426 0 126482 800
rect 129922 0 129978 800
rect 133326 0 133382 800
rect 136822 0 136878 800
rect 140318 0 140374 800
rect 143722 0 143778 800
rect 147218 0 147274 800
rect 150714 0 150770 800
rect 154118 0 154174 800
rect 157614 0 157670 800
rect 161110 0 161166 800
rect 164514 0 164570 800
rect 168010 0 168066 800
rect 171506 0 171562 800
rect 175002 0 175058 800
rect 178406 0 178462 800
rect 181902 0 181958 800
rect 185398 0 185454 800
rect 188802 0 188858 800
rect 192298 0 192354 800
rect 195794 0 195850 800
rect 199198 0 199254 800
rect 202694 0 202750 800
rect 206190 0 206246 800
rect 209594 0 209650 800
rect 213090 0 213146 800
rect 216586 0 216642 800
rect 219990 0 220046 800
rect 223486 0 223542 800
rect 226982 0 227038 800
rect 230386 0 230442 800
rect 233882 0 233938 800
rect 237378 0 237434 800
rect 240782 0 240838 800
rect 244278 0 244334 800
rect 247774 0 247830 800
rect 251178 0 251234 800
rect 254674 0 254730 800
rect 258170 0 258226 800
<< obsm2 >>
rect 572 856 258224 259593
rect 572 439 1618 856
rect 1786 439 5022 856
rect 5190 439 8518 856
rect 8686 439 12014 856
rect 12182 439 15418 856
rect 15586 439 18914 856
rect 19082 439 22410 856
rect 22578 439 25814 856
rect 25982 439 29310 856
rect 29478 439 32806 856
rect 32974 439 36210 856
rect 36378 439 39706 856
rect 39874 439 43202 856
rect 43370 439 46606 856
rect 46774 439 50102 856
rect 50270 439 53598 856
rect 53766 439 57002 856
rect 57170 439 60498 856
rect 60666 439 63994 856
rect 64162 439 67398 856
rect 67566 439 70894 856
rect 71062 439 74390 856
rect 74558 439 77794 856
rect 77962 439 81290 856
rect 81458 439 84786 856
rect 84954 439 88282 856
rect 88450 439 91686 856
rect 91854 439 95182 856
rect 95350 439 98678 856
rect 98846 439 102082 856
rect 102250 439 105578 856
rect 105746 439 109074 856
rect 109242 439 112478 856
rect 112646 439 115974 856
rect 116142 439 119470 856
rect 119638 439 122874 856
rect 123042 439 126370 856
rect 126538 439 129866 856
rect 130034 439 133270 856
rect 133438 439 136766 856
rect 136934 439 140262 856
rect 140430 439 143666 856
rect 143834 439 147162 856
rect 147330 439 150658 856
rect 150826 439 154062 856
rect 154230 439 157558 856
rect 157726 439 161054 856
rect 161222 439 164458 856
rect 164626 439 167954 856
rect 168122 439 171450 856
rect 171618 439 174946 856
rect 175114 439 178350 856
rect 178518 439 181846 856
rect 182014 439 185342 856
rect 185510 439 188746 856
rect 188914 439 192242 856
rect 192410 439 195738 856
rect 195906 439 199142 856
rect 199310 439 202638 856
rect 202806 439 206134 856
rect 206302 439 209538 856
rect 209706 439 213034 856
rect 213202 439 216530 856
rect 216698 439 219934 856
rect 220102 439 223430 856
rect 223598 439 226926 856
rect 227094 439 230330 856
rect 230498 439 233826 856
rect 233994 439 237322 856
rect 237490 439 240726 856
rect 240894 439 244222 856
rect 244390 439 247718 856
rect 247886 439 251122 856
rect 251290 439 254618 856
rect 254786 439 258114 856
<< metal3 >>
rect 0 259496 800 259616
rect 0 258680 800 258800
rect 0 257728 800 257848
rect 0 256912 800 257032
rect 0 255960 800 256080
rect 0 255144 800 255264
rect 0 254192 800 254312
rect 0 253376 800 253496
rect 0 252424 800 252544
rect 0 251608 800 251728
rect 0 250656 800 250776
rect 0 249840 800 249960
rect 0 249024 800 249144
rect 0 248072 800 248192
rect 0 247256 800 247376
rect 0 246304 800 246424
rect 0 245488 800 245608
rect 0 244536 800 244656
rect 0 243720 800 243840
rect 0 242768 800 242888
rect 0 241952 800 242072
rect 0 241000 800 241120
rect 0 240184 800 240304
rect 0 239232 800 239352
rect 0 238416 800 238536
rect 0 237600 800 237720
rect 0 236648 800 236768
rect 0 235832 800 235952
rect 0 234880 800 235000
rect 0 234064 800 234184
rect 0 233112 800 233232
rect 0 232296 800 232416
rect 0 231344 800 231464
rect 0 230528 800 230648
rect 0 229576 800 229696
rect 0 228760 800 228880
rect 0 227944 800 228064
rect 0 226992 800 227112
rect 0 226176 800 226296
rect 0 225224 800 225344
rect 0 224408 800 224528
rect 0 223456 800 223576
rect 0 222640 800 222760
rect 0 221688 800 221808
rect 0 220872 800 220992
rect 0 219920 800 220040
rect 0 219104 800 219224
rect 0 218152 800 218272
rect 0 217336 800 217456
rect 0 216520 800 216640
rect 0 215568 800 215688
rect 0 214752 800 214872
rect 0 213800 800 213920
rect 0 212984 800 213104
rect 0 212032 800 212152
rect 0 211216 800 211336
rect 0 210264 800 210384
rect 0 209448 800 209568
rect 0 208496 800 208616
rect 0 207680 800 207800
rect 0 206728 800 206848
rect 0 205912 800 206032
rect 0 205096 800 205216
rect 0 204144 800 204264
rect 0 203328 800 203448
rect 0 202376 800 202496
rect 0 201560 800 201680
rect 0 200608 800 200728
rect 0 199792 800 199912
rect 0 198840 800 198960
rect 0 198024 800 198144
rect 0 197072 800 197192
rect 0 196256 800 196376
rect 0 195440 800 195560
rect 0 194488 800 194608
rect 0 193672 800 193792
rect 0 192720 800 192840
rect 0 191904 800 192024
rect 0 190952 800 191072
rect 0 190136 800 190256
rect 0 189184 800 189304
rect 0 188368 800 188488
rect 0 187416 800 187536
rect 0 186600 800 186720
rect 0 185648 800 185768
rect 0 184832 800 184952
rect 0 184016 800 184136
rect 0 183064 800 183184
rect 0 182248 800 182368
rect 0 181296 800 181416
rect 0 180480 800 180600
rect 0 179528 800 179648
rect 0 178712 800 178832
rect 0 177760 800 177880
rect 0 176944 800 177064
rect 0 175992 800 176112
rect 0 175176 800 175296
rect 0 174224 800 174344
rect 0 173408 800 173528
rect 0 172592 800 172712
rect 0 171640 800 171760
rect 0 170824 800 170944
rect 0 169872 800 169992
rect 0 169056 800 169176
rect 0 168104 800 168224
rect 0 167288 800 167408
rect 0 166336 800 166456
rect 0 165520 800 165640
rect 0 164568 800 164688
rect 0 163752 800 163872
rect 0 162936 800 163056
rect 0 161984 800 162104
rect 0 161168 800 161288
rect 0 160216 800 160336
rect 0 159400 800 159520
rect 0 158448 800 158568
rect 0 157632 800 157752
rect 0 156680 800 156800
rect 0 155864 800 155984
rect 0 154912 800 155032
rect 0 154096 800 154216
rect 0 153144 800 153264
rect 0 152328 800 152448
rect 0 151512 800 151632
rect 0 150560 800 150680
rect 0 149744 800 149864
rect 0 148792 800 148912
rect 0 147976 800 148096
rect 0 147024 800 147144
rect 0 146208 800 146328
rect 0 145256 800 145376
rect 0 144440 800 144560
rect 0 143488 800 143608
rect 0 142672 800 142792
rect 0 141720 800 141840
rect 0 140904 800 141024
rect 0 140088 800 140208
rect 0 139136 800 139256
rect 0 138320 800 138440
rect 0 137368 800 137488
rect 0 136552 800 136672
rect 0 135600 800 135720
rect 0 134784 800 134904
rect 0 133832 800 133952
rect 0 133016 800 133136
rect 0 132064 800 132184
rect 0 131248 800 131368
rect 0 130432 800 130552
rect 0 129480 800 129600
rect 0 128664 800 128784
rect 0 127712 800 127832
rect 0 126896 800 127016
rect 0 125944 800 126064
rect 0 125128 800 125248
rect 0 124176 800 124296
rect 0 123360 800 123480
rect 0 122408 800 122528
rect 0 121592 800 121712
rect 0 120640 800 120760
rect 0 119824 800 119944
rect 0 119008 800 119128
rect 0 118056 800 118176
rect 0 117240 800 117360
rect 0 116288 800 116408
rect 0 115472 800 115592
rect 0 114520 800 114640
rect 0 113704 800 113824
rect 0 112752 800 112872
rect 0 111936 800 112056
rect 0 110984 800 111104
rect 0 110168 800 110288
rect 0 109216 800 109336
rect 0 108400 800 108520
rect 0 107584 800 107704
rect 0 106632 800 106752
rect 0 105816 800 105936
rect 0 104864 800 104984
rect 0 104048 800 104168
rect 0 103096 800 103216
rect 0 102280 800 102400
rect 0 101328 800 101448
rect 0 100512 800 100632
rect 0 99560 800 99680
rect 0 98744 800 98864
rect 0 97928 800 98048
rect 0 96976 800 97096
rect 0 96160 800 96280
rect 0 95208 800 95328
rect 0 94392 800 94512
rect 0 93440 800 93560
rect 0 92624 800 92744
rect 0 91672 800 91792
rect 0 90856 800 90976
rect 0 89904 800 90024
rect 0 89088 800 89208
rect 0 88136 800 88256
rect 0 87320 800 87440
rect 0 86504 800 86624
rect 0 85552 800 85672
rect 0 84736 800 84856
rect 0 83784 800 83904
rect 0 82968 800 83088
rect 0 82016 800 82136
rect 0 81200 800 81320
rect 0 80248 800 80368
rect 0 79432 800 79552
rect 0 78480 800 78600
rect 0 77664 800 77784
rect 0 76712 800 76832
rect 0 75896 800 76016
rect 0 75080 800 75200
rect 0 74128 800 74248
rect 0 73312 800 73432
rect 0 72360 800 72480
rect 0 71544 800 71664
rect 0 70592 800 70712
rect 0 69776 800 69896
rect 0 68824 800 68944
rect 0 68008 800 68128
rect 0 67056 800 67176
rect 0 66240 800 66360
rect 0 65424 800 65544
rect 0 64472 800 64592
rect 0 63656 800 63776
rect 0 62704 800 62824
rect 0 61888 800 62008
rect 0 60936 800 61056
rect 0 60120 800 60240
rect 0 59168 800 59288
rect 0 58352 800 58472
rect 0 57400 800 57520
rect 0 56584 800 56704
rect 0 55632 800 55752
rect 0 54816 800 54936
rect 0 54000 800 54120
rect 0 53048 800 53168
rect 0 52232 800 52352
rect 0 51280 800 51400
rect 0 50464 800 50584
rect 0 49512 800 49632
rect 0 48696 800 48816
rect 0 47744 800 47864
rect 0 46928 800 47048
rect 0 45976 800 46096
rect 0 45160 800 45280
rect 0 44208 800 44328
rect 0 43392 800 43512
rect 0 42576 800 42696
rect 0 41624 800 41744
rect 0 40808 800 40928
rect 0 39856 800 39976
rect 0 39040 800 39160
rect 0 38088 800 38208
rect 0 37272 800 37392
rect 0 36320 800 36440
rect 0 35504 800 35624
rect 0 34552 800 34672
rect 0 33736 800 33856
rect 0 32920 800 33040
rect 0 31968 800 32088
rect 0 31152 800 31272
rect 0 30200 800 30320
rect 0 29384 800 29504
rect 0 28432 800 28552
rect 0 27616 800 27736
rect 0 26664 800 26784
rect 0 25848 800 25968
rect 0 24896 800 25016
rect 0 24080 800 24200
rect 0 23128 800 23248
rect 0 22312 800 22432
rect 0 21496 800 21616
rect 0 20544 800 20664
rect 0 19728 800 19848
rect 0 18776 800 18896
rect 0 17960 800 18080
rect 0 17008 800 17128
rect 0 16192 800 16312
rect 0 15240 800 15360
rect 0 14424 800 14544
rect 0 13472 800 13592
rect 0 12656 800 12776
rect 0 11704 800 11824
rect 0 10888 800 11008
rect 0 10072 800 10192
rect 0 9120 800 9240
rect 0 8304 800 8424
rect 0 7352 800 7472
rect 0 6536 800 6656
rect 0 5584 800 5704
rect 0 4768 800 4888
rect 0 3816 800 3936
rect 0 3000 800 3120
rect 0 2048 800 2168
rect 0 1232 800 1352
rect 0 416 800 536
<< obsm3 >>
rect 880 259416 250288 259589
rect 606 258880 250288 259416
rect 880 258600 250288 258880
rect 606 257928 250288 258600
rect 880 257648 250288 257928
rect 606 257112 250288 257648
rect 880 256832 250288 257112
rect 606 256160 250288 256832
rect 880 255880 250288 256160
rect 606 255344 250288 255880
rect 880 255064 250288 255344
rect 606 254392 250288 255064
rect 880 254112 250288 254392
rect 606 253576 250288 254112
rect 880 253296 250288 253576
rect 606 252624 250288 253296
rect 880 252344 250288 252624
rect 606 251808 250288 252344
rect 880 251528 250288 251808
rect 606 250856 250288 251528
rect 880 250576 250288 250856
rect 606 250040 250288 250576
rect 880 249760 250288 250040
rect 606 249224 250288 249760
rect 880 248944 250288 249224
rect 606 248272 250288 248944
rect 880 247992 250288 248272
rect 606 247456 250288 247992
rect 880 247176 250288 247456
rect 606 246504 250288 247176
rect 880 246224 250288 246504
rect 606 245688 250288 246224
rect 880 245408 250288 245688
rect 606 244736 250288 245408
rect 880 244456 250288 244736
rect 606 243920 250288 244456
rect 880 243640 250288 243920
rect 606 242968 250288 243640
rect 880 242688 250288 242968
rect 606 242152 250288 242688
rect 880 241872 250288 242152
rect 606 241200 250288 241872
rect 880 240920 250288 241200
rect 606 240384 250288 240920
rect 880 240104 250288 240384
rect 606 239432 250288 240104
rect 880 239152 250288 239432
rect 606 238616 250288 239152
rect 880 238336 250288 238616
rect 606 237800 250288 238336
rect 880 237520 250288 237800
rect 606 236848 250288 237520
rect 880 236568 250288 236848
rect 606 236032 250288 236568
rect 880 235752 250288 236032
rect 606 235080 250288 235752
rect 880 234800 250288 235080
rect 606 234264 250288 234800
rect 880 233984 250288 234264
rect 606 233312 250288 233984
rect 880 233032 250288 233312
rect 606 232496 250288 233032
rect 880 232216 250288 232496
rect 606 231544 250288 232216
rect 880 231264 250288 231544
rect 606 230728 250288 231264
rect 880 230448 250288 230728
rect 606 229776 250288 230448
rect 880 229496 250288 229776
rect 606 228960 250288 229496
rect 880 228680 250288 228960
rect 606 228144 250288 228680
rect 880 227864 250288 228144
rect 606 227192 250288 227864
rect 880 226912 250288 227192
rect 606 226376 250288 226912
rect 880 226096 250288 226376
rect 606 225424 250288 226096
rect 880 225144 250288 225424
rect 606 224608 250288 225144
rect 880 224328 250288 224608
rect 606 223656 250288 224328
rect 880 223376 250288 223656
rect 606 222840 250288 223376
rect 880 222560 250288 222840
rect 606 221888 250288 222560
rect 880 221608 250288 221888
rect 606 221072 250288 221608
rect 880 220792 250288 221072
rect 606 220120 250288 220792
rect 880 219840 250288 220120
rect 606 219304 250288 219840
rect 880 219024 250288 219304
rect 606 218352 250288 219024
rect 880 218072 250288 218352
rect 606 217536 250288 218072
rect 880 217256 250288 217536
rect 606 216720 250288 217256
rect 880 216440 250288 216720
rect 606 215768 250288 216440
rect 880 215488 250288 215768
rect 606 214952 250288 215488
rect 880 214672 250288 214952
rect 606 214000 250288 214672
rect 880 213720 250288 214000
rect 606 213184 250288 213720
rect 880 212904 250288 213184
rect 606 212232 250288 212904
rect 880 211952 250288 212232
rect 606 211416 250288 211952
rect 880 211136 250288 211416
rect 606 210464 250288 211136
rect 880 210184 250288 210464
rect 606 209648 250288 210184
rect 880 209368 250288 209648
rect 606 208696 250288 209368
rect 880 208416 250288 208696
rect 606 207880 250288 208416
rect 880 207600 250288 207880
rect 606 206928 250288 207600
rect 880 206648 250288 206928
rect 606 206112 250288 206648
rect 880 205832 250288 206112
rect 606 205296 250288 205832
rect 880 205016 250288 205296
rect 606 204344 250288 205016
rect 880 204064 250288 204344
rect 606 203528 250288 204064
rect 880 203248 250288 203528
rect 606 202576 250288 203248
rect 880 202296 250288 202576
rect 606 201760 250288 202296
rect 880 201480 250288 201760
rect 606 200808 250288 201480
rect 880 200528 250288 200808
rect 606 199992 250288 200528
rect 880 199712 250288 199992
rect 606 199040 250288 199712
rect 880 198760 250288 199040
rect 606 198224 250288 198760
rect 880 197944 250288 198224
rect 606 197272 250288 197944
rect 880 196992 250288 197272
rect 606 196456 250288 196992
rect 880 196176 250288 196456
rect 606 195640 250288 196176
rect 880 195360 250288 195640
rect 606 194688 250288 195360
rect 880 194408 250288 194688
rect 606 193872 250288 194408
rect 880 193592 250288 193872
rect 606 192920 250288 193592
rect 880 192640 250288 192920
rect 606 192104 250288 192640
rect 880 191824 250288 192104
rect 606 191152 250288 191824
rect 880 190872 250288 191152
rect 606 190336 250288 190872
rect 880 190056 250288 190336
rect 606 189384 250288 190056
rect 880 189104 250288 189384
rect 606 188568 250288 189104
rect 880 188288 250288 188568
rect 606 187616 250288 188288
rect 880 187336 250288 187616
rect 606 186800 250288 187336
rect 880 186520 250288 186800
rect 606 185848 250288 186520
rect 880 185568 250288 185848
rect 606 185032 250288 185568
rect 880 184752 250288 185032
rect 606 184216 250288 184752
rect 880 183936 250288 184216
rect 606 183264 250288 183936
rect 880 182984 250288 183264
rect 606 182448 250288 182984
rect 880 182168 250288 182448
rect 606 181496 250288 182168
rect 880 181216 250288 181496
rect 606 180680 250288 181216
rect 880 180400 250288 180680
rect 606 179728 250288 180400
rect 880 179448 250288 179728
rect 606 178912 250288 179448
rect 880 178632 250288 178912
rect 606 177960 250288 178632
rect 880 177680 250288 177960
rect 606 177144 250288 177680
rect 880 176864 250288 177144
rect 606 176192 250288 176864
rect 880 175912 250288 176192
rect 606 175376 250288 175912
rect 880 175096 250288 175376
rect 606 174424 250288 175096
rect 880 174144 250288 174424
rect 606 173608 250288 174144
rect 880 173328 250288 173608
rect 606 172792 250288 173328
rect 880 172512 250288 172792
rect 606 171840 250288 172512
rect 880 171560 250288 171840
rect 606 171024 250288 171560
rect 880 170744 250288 171024
rect 606 170072 250288 170744
rect 880 169792 250288 170072
rect 606 169256 250288 169792
rect 880 168976 250288 169256
rect 606 168304 250288 168976
rect 880 168024 250288 168304
rect 606 167488 250288 168024
rect 880 167208 250288 167488
rect 606 166536 250288 167208
rect 880 166256 250288 166536
rect 606 165720 250288 166256
rect 880 165440 250288 165720
rect 606 164768 250288 165440
rect 880 164488 250288 164768
rect 606 163952 250288 164488
rect 880 163672 250288 163952
rect 606 163136 250288 163672
rect 880 162856 250288 163136
rect 606 162184 250288 162856
rect 880 161904 250288 162184
rect 606 161368 250288 161904
rect 880 161088 250288 161368
rect 606 160416 250288 161088
rect 880 160136 250288 160416
rect 606 159600 250288 160136
rect 880 159320 250288 159600
rect 606 158648 250288 159320
rect 880 158368 250288 158648
rect 606 157832 250288 158368
rect 880 157552 250288 157832
rect 606 156880 250288 157552
rect 880 156600 250288 156880
rect 606 156064 250288 156600
rect 880 155784 250288 156064
rect 606 155112 250288 155784
rect 880 154832 250288 155112
rect 606 154296 250288 154832
rect 880 154016 250288 154296
rect 606 153344 250288 154016
rect 880 153064 250288 153344
rect 606 152528 250288 153064
rect 880 152248 250288 152528
rect 606 151712 250288 152248
rect 880 151432 250288 151712
rect 606 150760 250288 151432
rect 880 150480 250288 150760
rect 606 149944 250288 150480
rect 880 149664 250288 149944
rect 606 148992 250288 149664
rect 880 148712 250288 148992
rect 606 148176 250288 148712
rect 880 147896 250288 148176
rect 606 147224 250288 147896
rect 880 146944 250288 147224
rect 606 146408 250288 146944
rect 880 146128 250288 146408
rect 606 145456 250288 146128
rect 880 145176 250288 145456
rect 606 144640 250288 145176
rect 880 144360 250288 144640
rect 606 143688 250288 144360
rect 880 143408 250288 143688
rect 606 142872 250288 143408
rect 880 142592 250288 142872
rect 606 141920 250288 142592
rect 880 141640 250288 141920
rect 606 141104 250288 141640
rect 880 140824 250288 141104
rect 606 140288 250288 140824
rect 880 140008 250288 140288
rect 606 139336 250288 140008
rect 880 139056 250288 139336
rect 606 138520 250288 139056
rect 880 138240 250288 138520
rect 606 137568 250288 138240
rect 880 137288 250288 137568
rect 606 136752 250288 137288
rect 880 136472 250288 136752
rect 606 135800 250288 136472
rect 880 135520 250288 135800
rect 606 134984 250288 135520
rect 880 134704 250288 134984
rect 606 134032 250288 134704
rect 880 133752 250288 134032
rect 606 133216 250288 133752
rect 880 132936 250288 133216
rect 606 132264 250288 132936
rect 880 131984 250288 132264
rect 606 131448 250288 131984
rect 880 131168 250288 131448
rect 606 130632 250288 131168
rect 880 130352 250288 130632
rect 606 129680 250288 130352
rect 880 129400 250288 129680
rect 606 128864 250288 129400
rect 880 128584 250288 128864
rect 606 127912 250288 128584
rect 880 127632 250288 127912
rect 606 127096 250288 127632
rect 880 126816 250288 127096
rect 606 126144 250288 126816
rect 880 125864 250288 126144
rect 606 125328 250288 125864
rect 880 125048 250288 125328
rect 606 124376 250288 125048
rect 880 124096 250288 124376
rect 606 123560 250288 124096
rect 880 123280 250288 123560
rect 606 122608 250288 123280
rect 880 122328 250288 122608
rect 606 121792 250288 122328
rect 880 121512 250288 121792
rect 606 120840 250288 121512
rect 880 120560 250288 120840
rect 606 120024 250288 120560
rect 880 119744 250288 120024
rect 606 119208 250288 119744
rect 880 118928 250288 119208
rect 606 118256 250288 118928
rect 880 117976 250288 118256
rect 606 117440 250288 117976
rect 880 117160 250288 117440
rect 606 116488 250288 117160
rect 880 116208 250288 116488
rect 606 115672 250288 116208
rect 880 115392 250288 115672
rect 606 114720 250288 115392
rect 880 114440 250288 114720
rect 606 113904 250288 114440
rect 880 113624 250288 113904
rect 606 112952 250288 113624
rect 880 112672 250288 112952
rect 606 112136 250288 112672
rect 880 111856 250288 112136
rect 606 111184 250288 111856
rect 880 110904 250288 111184
rect 606 110368 250288 110904
rect 880 110088 250288 110368
rect 606 109416 250288 110088
rect 880 109136 250288 109416
rect 606 108600 250288 109136
rect 880 108320 250288 108600
rect 606 107784 250288 108320
rect 880 107504 250288 107784
rect 606 106832 250288 107504
rect 880 106552 250288 106832
rect 606 106016 250288 106552
rect 880 105736 250288 106016
rect 606 105064 250288 105736
rect 880 104784 250288 105064
rect 606 104248 250288 104784
rect 880 103968 250288 104248
rect 606 103296 250288 103968
rect 880 103016 250288 103296
rect 606 102480 250288 103016
rect 880 102200 250288 102480
rect 606 101528 250288 102200
rect 880 101248 250288 101528
rect 606 100712 250288 101248
rect 880 100432 250288 100712
rect 606 99760 250288 100432
rect 880 99480 250288 99760
rect 606 98944 250288 99480
rect 880 98664 250288 98944
rect 606 98128 250288 98664
rect 880 97848 250288 98128
rect 606 97176 250288 97848
rect 880 96896 250288 97176
rect 606 96360 250288 96896
rect 880 96080 250288 96360
rect 606 95408 250288 96080
rect 880 95128 250288 95408
rect 606 94592 250288 95128
rect 880 94312 250288 94592
rect 606 93640 250288 94312
rect 880 93360 250288 93640
rect 606 92824 250288 93360
rect 880 92544 250288 92824
rect 606 91872 250288 92544
rect 880 91592 250288 91872
rect 606 91056 250288 91592
rect 880 90776 250288 91056
rect 606 90104 250288 90776
rect 880 89824 250288 90104
rect 606 89288 250288 89824
rect 880 89008 250288 89288
rect 606 88336 250288 89008
rect 880 88056 250288 88336
rect 606 87520 250288 88056
rect 880 87240 250288 87520
rect 606 86704 250288 87240
rect 880 86424 250288 86704
rect 606 85752 250288 86424
rect 880 85472 250288 85752
rect 606 84936 250288 85472
rect 880 84656 250288 84936
rect 606 83984 250288 84656
rect 880 83704 250288 83984
rect 606 83168 250288 83704
rect 880 82888 250288 83168
rect 606 82216 250288 82888
rect 880 81936 250288 82216
rect 606 81400 250288 81936
rect 880 81120 250288 81400
rect 606 80448 250288 81120
rect 880 80168 250288 80448
rect 606 79632 250288 80168
rect 880 79352 250288 79632
rect 606 78680 250288 79352
rect 880 78400 250288 78680
rect 606 77864 250288 78400
rect 880 77584 250288 77864
rect 606 76912 250288 77584
rect 880 76632 250288 76912
rect 606 76096 250288 76632
rect 880 75816 250288 76096
rect 606 75280 250288 75816
rect 880 75000 250288 75280
rect 606 74328 250288 75000
rect 880 74048 250288 74328
rect 606 73512 250288 74048
rect 880 73232 250288 73512
rect 606 72560 250288 73232
rect 880 72280 250288 72560
rect 606 71744 250288 72280
rect 880 71464 250288 71744
rect 606 70792 250288 71464
rect 880 70512 250288 70792
rect 606 69976 250288 70512
rect 880 69696 250288 69976
rect 606 69024 250288 69696
rect 880 68744 250288 69024
rect 606 68208 250288 68744
rect 880 67928 250288 68208
rect 606 67256 250288 67928
rect 880 66976 250288 67256
rect 606 66440 250288 66976
rect 880 66160 250288 66440
rect 606 65624 250288 66160
rect 880 65344 250288 65624
rect 606 64672 250288 65344
rect 880 64392 250288 64672
rect 606 63856 250288 64392
rect 880 63576 250288 63856
rect 606 62904 250288 63576
rect 880 62624 250288 62904
rect 606 62088 250288 62624
rect 880 61808 250288 62088
rect 606 61136 250288 61808
rect 880 60856 250288 61136
rect 606 60320 250288 60856
rect 880 60040 250288 60320
rect 606 59368 250288 60040
rect 880 59088 250288 59368
rect 606 58552 250288 59088
rect 880 58272 250288 58552
rect 606 57600 250288 58272
rect 880 57320 250288 57600
rect 606 56784 250288 57320
rect 880 56504 250288 56784
rect 606 55832 250288 56504
rect 880 55552 250288 55832
rect 606 55016 250288 55552
rect 880 54736 250288 55016
rect 606 54200 250288 54736
rect 880 53920 250288 54200
rect 606 53248 250288 53920
rect 880 52968 250288 53248
rect 606 52432 250288 52968
rect 880 52152 250288 52432
rect 606 51480 250288 52152
rect 880 51200 250288 51480
rect 606 50664 250288 51200
rect 880 50384 250288 50664
rect 606 49712 250288 50384
rect 880 49432 250288 49712
rect 606 48896 250288 49432
rect 880 48616 250288 48896
rect 606 47944 250288 48616
rect 880 47664 250288 47944
rect 606 47128 250288 47664
rect 880 46848 250288 47128
rect 606 46176 250288 46848
rect 880 45896 250288 46176
rect 606 45360 250288 45896
rect 880 45080 250288 45360
rect 606 44408 250288 45080
rect 880 44128 250288 44408
rect 606 43592 250288 44128
rect 880 43312 250288 43592
rect 606 42776 250288 43312
rect 880 42496 250288 42776
rect 606 41824 250288 42496
rect 880 41544 250288 41824
rect 606 41008 250288 41544
rect 880 40728 250288 41008
rect 606 40056 250288 40728
rect 880 39776 250288 40056
rect 606 39240 250288 39776
rect 880 38960 250288 39240
rect 606 38288 250288 38960
rect 880 38008 250288 38288
rect 606 37472 250288 38008
rect 880 37192 250288 37472
rect 606 36520 250288 37192
rect 880 36240 250288 36520
rect 606 35704 250288 36240
rect 880 35424 250288 35704
rect 606 34752 250288 35424
rect 880 34472 250288 34752
rect 606 33936 250288 34472
rect 880 33656 250288 33936
rect 606 33120 250288 33656
rect 880 32840 250288 33120
rect 606 32168 250288 32840
rect 880 31888 250288 32168
rect 606 31352 250288 31888
rect 880 31072 250288 31352
rect 606 30400 250288 31072
rect 880 30120 250288 30400
rect 606 29584 250288 30120
rect 880 29304 250288 29584
rect 606 28632 250288 29304
rect 880 28352 250288 28632
rect 606 27816 250288 28352
rect 880 27536 250288 27816
rect 606 26864 250288 27536
rect 880 26584 250288 26864
rect 606 26048 250288 26584
rect 880 25768 250288 26048
rect 606 25096 250288 25768
rect 880 24816 250288 25096
rect 606 24280 250288 24816
rect 880 24000 250288 24280
rect 606 23328 250288 24000
rect 880 23048 250288 23328
rect 606 22512 250288 23048
rect 880 22232 250288 22512
rect 606 21696 250288 22232
rect 880 21416 250288 21696
rect 606 20744 250288 21416
rect 880 20464 250288 20744
rect 606 19928 250288 20464
rect 880 19648 250288 19928
rect 606 18976 250288 19648
rect 880 18696 250288 18976
rect 606 18160 250288 18696
rect 880 17880 250288 18160
rect 606 17208 250288 17880
rect 880 16928 250288 17208
rect 606 16392 250288 16928
rect 880 16112 250288 16392
rect 606 15440 250288 16112
rect 880 15160 250288 15440
rect 606 14624 250288 15160
rect 880 14344 250288 14624
rect 606 13672 250288 14344
rect 880 13392 250288 13672
rect 606 12856 250288 13392
rect 880 12576 250288 12856
rect 606 11904 250288 12576
rect 880 11624 250288 11904
rect 606 11088 250288 11624
rect 880 10808 250288 11088
rect 606 10272 250288 10808
rect 880 9992 250288 10272
rect 606 9320 250288 9992
rect 880 9040 250288 9320
rect 606 8504 250288 9040
rect 880 8224 250288 8504
rect 606 7552 250288 8224
rect 880 7272 250288 7552
rect 606 6736 250288 7272
rect 880 6456 250288 6736
rect 606 5784 250288 6456
rect 880 5504 250288 5784
rect 606 4968 250288 5504
rect 880 4688 250288 4968
rect 606 4016 250288 4688
rect 880 3736 250288 4016
rect 606 3200 250288 3736
rect 880 2920 250288 3200
rect 606 2248 250288 2920
rect 880 1968 250288 2248
rect 606 1432 250288 1968
rect 880 1152 250288 1432
rect 606 616 250288 1152
rect 880 443 250288 616
<< metal4 >>
rect 4208 2128 4528 257360
rect 19568 2128 19888 257360
rect 34928 2128 35248 257360
rect 50288 2128 50608 257360
rect 65648 2128 65968 257360
rect 81008 2128 81328 257360
rect 96368 2128 96688 257360
rect 111728 2128 112048 257360
rect 127088 2128 127408 257360
rect 142448 2128 142768 257360
rect 157808 2128 158128 257360
rect 173168 2128 173488 257360
rect 188528 2128 188848 257360
rect 203888 2128 204208 257360
rect 219248 2128 219568 257360
rect 234608 2128 234928 257360
rect 249968 2128 250288 257360
<< obsm4 >>
rect 611 2347 4128 254693
rect 4608 2347 19488 254693
rect 19968 2347 34848 254693
rect 35328 2347 50208 254693
rect 50688 2347 65568 254693
rect 66048 2347 80928 254693
rect 81408 2347 96288 254693
rect 96768 2347 111648 254693
rect 112128 2347 127008 254693
rect 127488 2347 142368 254693
rect 142848 2347 157728 254693
rect 158208 2347 173088 254693
rect 173568 2347 188448 254693
rect 188928 2347 202709 254693
<< labels >>
rlabel metal3 s 0 116288 800 116408 6 bb_addr0[0]
port 1 nsew signal output
rlabel metal3 s 0 163752 800 163872 6 bb_addr0[10]
port 2 nsew signal output
rlabel metal3 s 0 168104 800 168224 6 bb_addr0[11]
port 3 nsew signal output
rlabel metal3 s 0 172592 800 172712 6 bb_addr0[12]
port 4 nsew signal output
rlabel metal3 s 0 176944 800 177064 6 bb_addr0[13]
port 5 nsew signal output
rlabel metal3 s 0 181296 800 181416 6 bb_addr0[14]
port 6 nsew signal output
rlabel metal3 s 0 185648 800 185768 6 bb_addr0[15]
port 7 nsew signal output
rlabel metal3 s 0 190136 800 190256 6 bb_addr0[16]
port 8 nsew signal output
rlabel metal3 s 0 194488 800 194608 6 bb_addr0[17]
port 9 nsew signal output
rlabel metal3 s 0 198840 800 198960 6 bb_addr0[18]
port 10 nsew signal output
rlabel metal3 s 0 203328 800 203448 6 bb_addr0[19]
port 11 nsew signal output
rlabel metal3 s 0 121592 800 121712 6 bb_addr0[1]
port 12 nsew signal output
rlabel metal3 s 0 207680 800 207800 6 bb_addr0[20]
port 13 nsew signal output
rlabel metal3 s 0 212032 800 212152 6 bb_addr0[21]
port 14 nsew signal output
rlabel metal3 s 0 216520 800 216640 6 bb_addr0[22]
port 15 nsew signal output
rlabel metal3 s 0 220872 800 220992 6 bb_addr0[23]
port 16 nsew signal output
rlabel metal3 s 0 225224 800 225344 6 bb_addr0[24]
port 17 nsew signal output
rlabel metal3 s 0 229576 800 229696 6 bb_addr0[25]
port 18 nsew signal output
rlabel metal3 s 0 234064 800 234184 6 bb_addr0[26]
port 19 nsew signal output
rlabel metal3 s 0 238416 800 238536 6 bb_addr0[27]
port 20 nsew signal output
rlabel metal3 s 0 242768 800 242888 6 bb_addr0[28]
port 21 nsew signal output
rlabel metal3 s 0 247256 800 247376 6 bb_addr0[29]
port 22 nsew signal output
rlabel metal3 s 0 126896 800 127016 6 bb_addr0[2]
port 23 nsew signal output
rlabel metal3 s 0 251608 800 251728 6 bb_addr0[30]
port 24 nsew signal output
rlabel metal3 s 0 255960 800 256080 6 bb_addr0[31]
port 25 nsew signal output
rlabel metal3 s 0 132064 800 132184 6 bb_addr0[3]
port 26 nsew signal output
rlabel metal3 s 0 137368 800 137488 6 bb_addr0[4]
port 27 nsew signal output
rlabel metal3 s 0 141720 800 141840 6 bb_addr0[5]
port 28 nsew signal output
rlabel metal3 s 0 146208 800 146328 6 bb_addr0[6]
port 29 nsew signal output
rlabel metal3 s 0 150560 800 150680 6 bb_addr0[7]
port 30 nsew signal output
rlabel metal3 s 0 154912 800 155032 6 bb_addr0[8]
port 31 nsew signal output
rlabel metal3 s 0 159400 800 159520 6 bb_addr0[9]
port 32 nsew signal output
rlabel metal3 s 0 117240 800 117360 6 bb_addr1[0]
port 33 nsew signal output
rlabel metal3 s 0 164568 800 164688 6 bb_addr1[10]
port 34 nsew signal output
rlabel metal3 s 0 169056 800 169176 6 bb_addr1[11]
port 35 nsew signal output
rlabel metal3 s 0 173408 800 173528 6 bb_addr1[12]
port 36 nsew signal output
rlabel metal3 s 0 177760 800 177880 6 bb_addr1[13]
port 37 nsew signal output
rlabel metal3 s 0 182248 800 182368 6 bb_addr1[14]
port 38 nsew signal output
rlabel metal3 s 0 186600 800 186720 6 bb_addr1[15]
port 39 nsew signal output
rlabel metal3 s 0 190952 800 191072 6 bb_addr1[16]
port 40 nsew signal output
rlabel metal3 s 0 195440 800 195560 6 bb_addr1[17]
port 41 nsew signal output
rlabel metal3 s 0 199792 800 199912 6 bb_addr1[18]
port 42 nsew signal output
rlabel metal3 s 0 204144 800 204264 6 bb_addr1[19]
port 43 nsew signal output
rlabel metal3 s 0 122408 800 122528 6 bb_addr1[1]
port 44 nsew signal output
rlabel metal3 s 0 208496 800 208616 6 bb_addr1[20]
port 45 nsew signal output
rlabel metal3 s 0 212984 800 213104 6 bb_addr1[21]
port 46 nsew signal output
rlabel metal3 s 0 217336 800 217456 6 bb_addr1[22]
port 47 nsew signal output
rlabel metal3 s 0 221688 800 221808 6 bb_addr1[23]
port 48 nsew signal output
rlabel metal3 s 0 226176 800 226296 6 bb_addr1[24]
port 49 nsew signal output
rlabel metal3 s 0 230528 800 230648 6 bb_addr1[25]
port 50 nsew signal output
rlabel metal3 s 0 234880 800 235000 6 bb_addr1[26]
port 51 nsew signal output
rlabel metal3 s 0 239232 800 239352 6 bb_addr1[27]
port 52 nsew signal output
rlabel metal3 s 0 243720 800 243840 6 bb_addr1[28]
port 53 nsew signal output
rlabel metal3 s 0 248072 800 248192 6 bb_addr1[29]
port 54 nsew signal output
rlabel metal3 s 0 127712 800 127832 6 bb_addr1[2]
port 55 nsew signal output
rlabel metal3 s 0 252424 800 252544 6 bb_addr1[30]
port 56 nsew signal output
rlabel metal3 s 0 256912 800 257032 6 bb_addr1[31]
port 57 nsew signal output
rlabel metal3 s 0 133016 800 133136 6 bb_addr1[3]
port 58 nsew signal output
rlabel metal3 s 0 138320 800 138440 6 bb_addr1[4]
port 59 nsew signal output
rlabel metal3 s 0 142672 800 142792 6 bb_addr1[5]
port 60 nsew signal output
rlabel metal3 s 0 147024 800 147144 6 bb_addr1[6]
port 61 nsew signal output
rlabel metal3 s 0 151512 800 151632 6 bb_addr1[7]
port 62 nsew signal output
rlabel metal3 s 0 155864 800 155984 6 bb_addr1[8]
port 63 nsew signal output
rlabel metal3 s 0 160216 800 160336 6 bb_addr1[9]
port 64 nsew signal output
rlabel metal3 s 0 113704 800 113824 6 bb_csb0
port 65 nsew signal output
rlabel metal3 s 0 114520 800 114640 6 bb_csb1
port 66 nsew signal output
rlabel metal3 s 0 118056 800 118176 6 bb_din0[0]
port 67 nsew signal output
rlabel metal3 s 0 165520 800 165640 6 bb_din0[10]
port 68 nsew signal output
rlabel metal3 s 0 169872 800 169992 6 bb_din0[11]
port 69 nsew signal output
rlabel metal3 s 0 174224 800 174344 6 bb_din0[12]
port 70 nsew signal output
rlabel metal3 s 0 178712 800 178832 6 bb_din0[13]
port 71 nsew signal output
rlabel metal3 s 0 183064 800 183184 6 bb_din0[14]
port 72 nsew signal output
rlabel metal3 s 0 187416 800 187536 6 bb_din0[15]
port 73 nsew signal output
rlabel metal3 s 0 191904 800 192024 6 bb_din0[16]
port 74 nsew signal output
rlabel metal3 s 0 196256 800 196376 6 bb_din0[17]
port 75 nsew signal output
rlabel metal3 s 0 200608 800 200728 6 bb_din0[18]
port 76 nsew signal output
rlabel metal3 s 0 205096 800 205216 6 bb_din0[19]
port 77 nsew signal output
rlabel metal3 s 0 123360 800 123480 6 bb_din0[1]
port 78 nsew signal output
rlabel metal3 s 0 209448 800 209568 6 bb_din0[20]
port 79 nsew signal output
rlabel metal3 s 0 213800 800 213920 6 bb_din0[21]
port 80 nsew signal output
rlabel metal3 s 0 218152 800 218272 6 bb_din0[22]
port 81 nsew signal output
rlabel metal3 s 0 222640 800 222760 6 bb_din0[23]
port 82 nsew signal output
rlabel metal3 s 0 226992 800 227112 6 bb_din0[24]
port 83 nsew signal output
rlabel metal3 s 0 231344 800 231464 6 bb_din0[25]
port 84 nsew signal output
rlabel metal3 s 0 235832 800 235952 6 bb_din0[26]
port 85 nsew signal output
rlabel metal3 s 0 240184 800 240304 6 bb_din0[27]
port 86 nsew signal output
rlabel metal3 s 0 244536 800 244656 6 bb_din0[28]
port 87 nsew signal output
rlabel metal3 s 0 249024 800 249144 6 bb_din0[29]
port 88 nsew signal output
rlabel metal3 s 0 128664 800 128784 6 bb_din0[2]
port 89 nsew signal output
rlabel metal3 s 0 253376 800 253496 6 bb_din0[30]
port 90 nsew signal output
rlabel metal3 s 0 257728 800 257848 6 bb_din0[31]
port 91 nsew signal output
rlabel metal3 s 0 133832 800 133952 6 bb_din0[3]
port 92 nsew signal output
rlabel metal3 s 0 139136 800 139256 6 bb_din0[4]
port 93 nsew signal output
rlabel metal3 s 0 143488 800 143608 6 bb_din0[5]
port 94 nsew signal output
rlabel metal3 s 0 147976 800 148096 6 bb_din0[6]
port 95 nsew signal output
rlabel metal3 s 0 152328 800 152448 6 bb_din0[7]
port 96 nsew signal output
rlabel metal3 s 0 156680 800 156800 6 bb_din0[8]
port 97 nsew signal output
rlabel metal3 s 0 161168 800 161288 6 bb_din0[9]
port 98 nsew signal output
rlabel metal3 s 0 119008 800 119128 6 bb_dout0[0]
port 99 nsew signal input
rlabel metal3 s 0 166336 800 166456 6 bb_dout0[10]
port 100 nsew signal input
rlabel metal3 s 0 170824 800 170944 6 bb_dout0[11]
port 101 nsew signal input
rlabel metal3 s 0 175176 800 175296 6 bb_dout0[12]
port 102 nsew signal input
rlabel metal3 s 0 179528 800 179648 6 bb_dout0[13]
port 103 nsew signal input
rlabel metal3 s 0 184016 800 184136 6 bb_dout0[14]
port 104 nsew signal input
rlabel metal3 s 0 188368 800 188488 6 bb_dout0[15]
port 105 nsew signal input
rlabel metal3 s 0 192720 800 192840 6 bb_dout0[16]
port 106 nsew signal input
rlabel metal3 s 0 197072 800 197192 6 bb_dout0[17]
port 107 nsew signal input
rlabel metal3 s 0 201560 800 201680 6 bb_dout0[18]
port 108 nsew signal input
rlabel metal3 s 0 205912 800 206032 6 bb_dout0[19]
port 109 nsew signal input
rlabel metal3 s 0 124176 800 124296 6 bb_dout0[1]
port 110 nsew signal input
rlabel metal3 s 0 210264 800 210384 6 bb_dout0[20]
port 111 nsew signal input
rlabel metal3 s 0 214752 800 214872 6 bb_dout0[21]
port 112 nsew signal input
rlabel metal3 s 0 219104 800 219224 6 bb_dout0[22]
port 113 nsew signal input
rlabel metal3 s 0 223456 800 223576 6 bb_dout0[23]
port 114 nsew signal input
rlabel metal3 s 0 227944 800 228064 6 bb_dout0[24]
port 115 nsew signal input
rlabel metal3 s 0 232296 800 232416 6 bb_dout0[25]
port 116 nsew signal input
rlabel metal3 s 0 236648 800 236768 6 bb_dout0[26]
port 117 nsew signal input
rlabel metal3 s 0 241000 800 241120 6 bb_dout0[27]
port 118 nsew signal input
rlabel metal3 s 0 245488 800 245608 6 bb_dout0[28]
port 119 nsew signal input
rlabel metal3 s 0 249840 800 249960 6 bb_dout0[29]
port 120 nsew signal input
rlabel metal3 s 0 129480 800 129600 6 bb_dout0[2]
port 121 nsew signal input
rlabel metal3 s 0 254192 800 254312 6 bb_dout0[30]
port 122 nsew signal input
rlabel metal3 s 0 258680 800 258800 6 bb_dout0[31]
port 123 nsew signal input
rlabel metal3 s 0 134784 800 134904 6 bb_dout0[3]
port 124 nsew signal input
rlabel metal3 s 0 140088 800 140208 6 bb_dout0[4]
port 125 nsew signal input
rlabel metal3 s 0 144440 800 144560 6 bb_dout0[5]
port 126 nsew signal input
rlabel metal3 s 0 148792 800 148912 6 bb_dout0[6]
port 127 nsew signal input
rlabel metal3 s 0 153144 800 153264 6 bb_dout0[7]
port 128 nsew signal input
rlabel metal3 s 0 157632 800 157752 6 bb_dout0[8]
port 129 nsew signal input
rlabel metal3 s 0 161984 800 162104 6 bb_dout0[9]
port 130 nsew signal input
rlabel metal3 s 0 119824 800 119944 6 bb_dout1[0]
port 131 nsew signal input
rlabel metal3 s 0 167288 800 167408 6 bb_dout1[10]
port 132 nsew signal input
rlabel metal3 s 0 171640 800 171760 6 bb_dout1[11]
port 133 nsew signal input
rlabel metal3 s 0 175992 800 176112 6 bb_dout1[12]
port 134 nsew signal input
rlabel metal3 s 0 180480 800 180600 6 bb_dout1[13]
port 135 nsew signal input
rlabel metal3 s 0 184832 800 184952 6 bb_dout1[14]
port 136 nsew signal input
rlabel metal3 s 0 189184 800 189304 6 bb_dout1[15]
port 137 nsew signal input
rlabel metal3 s 0 193672 800 193792 6 bb_dout1[16]
port 138 nsew signal input
rlabel metal3 s 0 198024 800 198144 6 bb_dout1[17]
port 139 nsew signal input
rlabel metal3 s 0 202376 800 202496 6 bb_dout1[18]
port 140 nsew signal input
rlabel metal3 s 0 206728 800 206848 6 bb_dout1[19]
port 141 nsew signal input
rlabel metal3 s 0 125128 800 125248 6 bb_dout1[1]
port 142 nsew signal input
rlabel metal3 s 0 211216 800 211336 6 bb_dout1[20]
port 143 nsew signal input
rlabel metal3 s 0 215568 800 215688 6 bb_dout1[21]
port 144 nsew signal input
rlabel metal3 s 0 219920 800 220040 6 bb_dout1[22]
port 145 nsew signal input
rlabel metal3 s 0 224408 800 224528 6 bb_dout1[23]
port 146 nsew signal input
rlabel metal3 s 0 228760 800 228880 6 bb_dout1[24]
port 147 nsew signal input
rlabel metal3 s 0 233112 800 233232 6 bb_dout1[25]
port 148 nsew signal input
rlabel metal3 s 0 237600 800 237720 6 bb_dout1[26]
port 149 nsew signal input
rlabel metal3 s 0 241952 800 242072 6 bb_dout1[27]
port 150 nsew signal input
rlabel metal3 s 0 246304 800 246424 6 bb_dout1[28]
port 151 nsew signal input
rlabel metal3 s 0 250656 800 250776 6 bb_dout1[29]
port 152 nsew signal input
rlabel metal3 s 0 130432 800 130552 6 bb_dout1[2]
port 153 nsew signal input
rlabel metal3 s 0 255144 800 255264 6 bb_dout1[30]
port 154 nsew signal input
rlabel metal3 s 0 259496 800 259616 6 bb_dout1[31]
port 155 nsew signal input
rlabel metal3 s 0 135600 800 135720 6 bb_dout1[3]
port 156 nsew signal input
rlabel metal3 s 0 140904 800 141024 6 bb_dout1[4]
port 157 nsew signal input
rlabel metal3 s 0 145256 800 145376 6 bb_dout1[5]
port 158 nsew signal input
rlabel metal3 s 0 149744 800 149864 6 bb_dout1[6]
port 159 nsew signal input
rlabel metal3 s 0 154096 800 154216 6 bb_dout1[7]
port 160 nsew signal input
rlabel metal3 s 0 158448 800 158568 6 bb_dout1[8]
port 161 nsew signal input
rlabel metal3 s 0 162936 800 163056 6 bb_dout1[9]
port 162 nsew signal input
rlabel metal3 s 0 115472 800 115592 6 bb_web0
port 163 nsew signal output
rlabel metal3 s 0 120640 800 120760 6 bb_wmask0[0]
port 164 nsew signal output
rlabel metal3 s 0 125944 800 126064 6 bb_wmask0[1]
port 165 nsew signal output
rlabel metal3 s 0 131248 800 131368 6 bb_wmask0[2]
port 166 nsew signal output
rlabel metal3 s 0 136552 800 136672 6 bb_wmask0[3]
port 167 nsew signal output
rlabel metal2 s 1674 0 1730 800 6 clk_g
port 168 nsew signal input
rlabel metal2 s 15474 0 15530 800 6 io_gecerli
port 169 nsew signal output
rlabel metal2 s 18970 0 19026 800 6 io_oeb[0]
port 170 nsew signal output
rlabel metal2 s 88338 0 88394 800 6 io_oeb[10]
port 171 nsew signal output
rlabel metal2 s 95238 0 95294 800 6 io_oeb[11]
port 172 nsew signal output
rlabel metal2 s 102138 0 102194 800 6 io_oeb[12]
port 173 nsew signal output
rlabel metal2 s 109130 0 109186 800 6 io_oeb[13]
port 174 nsew signal output
rlabel metal2 s 116030 0 116086 800 6 io_oeb[14]
port 175 nsew signal output
rlabel metal2 s 122930 0 122986 800 6 io_oeb[15]
port 176 nsew signal output
rlabel metal2 s 129922 0 129978 800 6 io_oeb[16]
port 177 nsew signal output
rlabel metal2 s 136822 0 136878 800 6 io_oeb[17]
port 178 nsew signal output
rlabel metal2 s 143722 0 143778 800 6 io_oeb[18]
port 179 nsew signal output
rlabel metal2 s 150714 0 150770 800 6 io_oeb[19]
port 180 nsew signal output
rlabel metal2 s 25870 0 25926 800 6 io_oeb[1]
port 181 nsew signal output
rlabel metal2 s 157614 0 157670 800 6 io_oeb[20]
port 182 nsew signal output
rlabel metal2 s 164514 0 164570 800 6 io_oeb[21]
port 183 nsew signal output
rlabel metal2 s 171506 0 171562 800 6 io_oeb[22]
port 184 nsew signal output
rlabel metal2 s 178406 0 178462 800 6 io_oeb[23]
port 185 nsew signal output
rlabel metal2 s 185398 0 185454 800 6 io_oeb[24]
port 186 nsew signal output
rlabel metal2 s 192298 0 192354 800 6 io_oeb[25]
port 187 nsew signal output
rlabel metal2 s 199198 0 199254 800 6 io_oeb[26]
port 188 nsew signal output
rlabel metal2 s 206190 0 206246 800 6 io_oeb[27]
port 189 nsew signal output
rlabel metal2 s 213090 0 213146 800 6 io_oeb[28]
port 190 nsew signal output
rlabel metal2 s 219990 0 220046 800 6 io_oeb[29]
port 191 nsew signal output
rlabel metal2 s 32862 0 32918 800 6 io_oeb[2]
port 192 nsew signal output
rlabel metal2 s 226982 0 227038 800 6 io_oeb[30]
port 193 nsew signal output
rlabel metal2 s 233882 0 233938 800 6 io_oeb[31]
port 194 nsew signal output
rlabel metal2 s 240782 0 240838 800 6 io_oeb[32]
port 195 nsew signal output
rlabel metal2 s 244278 0 244334 800 6 io_oeb[33]
port 196 nsew signal output
rlabel metal2 s 247774 0 247830 800 6 io_oeb[34]
port 197 nsew signal output
rlabel metal2 s 251178 0 251234 800 6 io_oeb[35]
port 198 nsew signal output
rlabel metal2 s 254674 0 254730 800 6 io_oeb[36]
port 199 nsew signal output
rlabel metal2 s 258170 0 258226 800 6 io_oeb[37]
port 200 nsew signal output
rlabel metal2 s 39762 0 39818 800 6 io_oeb[3]
port 201 nsew signal output
rlabel metal2 s 46662 0 46718 800 6 io_oeb[4]
port 202 nsew signal output
rlabel metal2 s 53654 0 53710 800 6 io_oeb[5]
port 203 nsew signal output
rlabel metal2 s 60554 0 60610 800 6 io_oeb[6]
port 204 nsew signal output
rlabel metal2 s 67454 0 67510 800 6 io_oeb[7]
port 205 nsew signal output
rlabel metal2 s 74446 0 74502 800 6 io_oeb[8]
port 206 nsew signal output
rlabel metal2 s 81346 0 81402 800 6 io_oeb[9]
port 207 nsew signal output
rlabel metal2 s 22466 0 22522 800 6 io_ps[0]
port 208 nsew signal output
rlabel metal2 s 91742 0 91798 800 6 io_ps[10]
port 209 nsew signal output
rlabel metal2 s 98734 0 98790 800 6 io_ps[11]
port 210 nsew signal output
rlabel metal2 s 105634 0 105690 800 6 io_ps[12]
port 211 nsew signal output
rlabel metal2 s 112534 0 112590 800 6 io_ps[13]
port 212 nsew signal output
rlabel metal2 s 119526 0 119582 800 6 io_ps[14]
port 213 nsew signal output
rlabel metal2 s 126426 0 126482 800 6 io_ps[15]
port 214 nsew signal output
rlabel metal2 s 133326 0 133382 800 6 io_ps[16]
port 215 nsew signal output
rlabel metal2 s 140318 0 140374 800 6 io_ps[17]
port 216 nsew signal output
rlabel metal2 s 147218 0 147274 800 6 io_ps[18]
port 217 nsew signal output
rlabel metal2 s 154118 0 154174 800 6 io_ps[19]
port 218 nsew signal output
rlabel metal2 s 29366 0 29422 800 6 io_ps[1]
port 219 nsew signal output
rlabel metal2 s 161110 0 161166 800 6 io_ps[20]
port 220 nsew signal output
rlabel metal2 s 168010 0 168066 800 6 io_ps[21]
port 221 nsew signal output
rlabel metal2 s 175002 0 175058 800 6 io_ps[22]
port 222 nsew signal output
rlabel metal2 s 181902 0 181958 800 6 io_ps[23]
port 223 nsew signal output
rlabel metal2 s 188802 0 188858 800 6 io_ps[24]
port 224 nsew signal output
rlabel metal2 s 195794 0 195850 800 6 io_ps[25]
port 225 nsew signal output
rlabel metal2 s 202694 0 202750 800 6 io_ps[26]
port 226 nsew signal output
rlabel metal2 s 209594 0 209650 800 6 io_ps[27]
port 227 nsew signal output
rlabel metal2 s 216586 0 216642 800 6 io_ps[28]
port 228 nsew signal output
rlabel metal2 s 223486 0 223542 800 6 io_ps[29]
port 229 nsew signal output
rlabel metal2 s 36266 0 36322 800 6 io_ps[2]
port 230 nsew signal output
rlabel metal2 s 230386 0 230442 800 6 io_ps[30]
port 231 nsew signal output
rlabel metal2 s 237378 0 237434 800 6 io_ps[31]
port 232 nsew signal output
rlabel metal2 s 43258 0 43314 800 6 io_ps[3]
port 233 nsew signal output
rlabel metal2 s 50158 0 50214 800 6 io_ps[4]
port 234 nsew signal output
rlabel metal2 s 57058 0 57114 800 6 io_ps[5]
port 235 nsew signal output
rlabel metal2 s 64050 0 64106 800 6 io_ps[6]
port 236 nsew signal output
rlabel metal2 s 70950 0 71006 800 6 io_ps[7]
port 237 nsew signal output
rlabel metal2 s 77850 0 77906 800 6 io_ps[8]
port 238 nsew signal output
rlabel metal2 s 84842 0 84898 800 6 io_ps[9]
port 239 nsew signal output
rlabel metal2 s 5078 0 5134 800 6 rst_g
port 240 nsew signal input
rlabel metal2 s 12070 0 12126 800 6 rx
port 241 nsew signal input
rlabel metal2 s 8574 0 8630 800 6 tx
port 242 nsew signal output
rlabel metal3 s 0 3000 800 3120 6 vb_addr0[0]
port 243 nsew signal output
rlabel metal3 s 0 50464 800 50584 6 vb_addr0[10]
port 244 nsew signal output
rlabel metal3 s 0 54816 800 54936 6 vb_addr0[11]
port 245 nsew signal output
rlabel metal3 s 0 59168 800 59288 6 vb_addr0[12]
port 246 nsew signal output
rlabel metal3 s 0 8304 800 8424 6 vb_addr0[1]
port 247 nsew signal output
rlabel metal3 s 0 13472 800 13592 6 vb_addr0[2]
port 248 nsew signal output
rlabel metal3 s 0 18776 800 18896 6 vb_addr0[3]
port 249 nsew signal output
rlabel metal3 s 0 24080 800 24200 6 vb_addr0[4]
port 250 nsew signal output
rlabel metal3 s 0 28432 800 28552 6 vb_addr0[5]
port 251 nsew signal output
rlabel metal3 s 0 32920 800 33040 6 vb_addr0[6]
port 252 nsew signal output
rlabel metal3 s 0 37272 800 37392 6 vb_addr0[7]
port 253 nsew signal output
rlabel metal3 s 0 41624 800 41744 6 vb_addr0[8]
port 254 nsew signal output
rlabel metal3 s 0 45976 800 46096 6 vb_addr0[9]
port 255 nsew signal output
rlabel metal3 s 0 3816 800 3936 6 vb_addr1[0]
port 256 nsew signal output
rlabel metal3 s 0 51280 800 51400 6 vb_addr1[10]
port 257 nsew signal output
rlabel metal3 s 0 55632 800 55752 6 vb_addr1[11]
port 258 nsew signal output
rlabel metal3 s 0 60120 800 60240 6 vb_addr1[12]
port 259 nsew signal output
rlabel metal3 s 0 9120 800 9240 6 vb_addr1[1]
port 260 nsew signal output
rlabel metal3 s 0 14424 800 14544 6 vb_addr1[2]
port 261 nsew signal output
rlabel metal3 s 0 19728 800 19848 6 vb_addr1[3]
port 262 nsew signal output
rlabel metal3 s 0 24896 800 25016 6 vb_addr1[4]
port 263 nsew signal output
rlabel metal3 s 0 29384 800 29504 6 vb_addr1[5]
port 264 nsew signal output
rlabel metal3 s 0 33736 800 33856 6 vb_addr1[6]
port 265 nsew signal output
rlabel metal3 s 0 38088 800 38208 6 vb_addr1[7]
port 266 nsew signal output
rlabel metal3 s 0 42576 800 42696 6 vb_addr1[8]
port 267 nsew signal output
rlabel metal3 s 0 46928 800 47048 6 vb_addr1[9]
port 268 nsew signal output
rlabel metal3 s 0 416 800 536 6 vb_csb0
port 269 nsew signal output
rlabel metal3 s 0 1232 800 1352 6 vb_csb1
port 270 nsew signal output
rlabel metal3 s 0 4768 800 4888 6 vb_din0[0]
port 271 nsew signal output
rlabel metal3 s 0 52232 800 52352 6 vb_din0[10]
port 272 nsew signal output
rlabel metal3 s 0 56584 800 56704 6 vb_din0[11]
port 273 nsew signal output
rlabel metal3 s 0 60936 800 61056 6 vb_din0[12]
port 274 nsew signal output
rlabel metal3 s 0 63656 800 63776 6 vb_din0[13]
port 275 nsew signal output
rlabel metal3 s 0 66240 800 66360 6 vb_din0[14]
port 276 nsew signal output
rlabel metal3 s 0 68824 800 68944 6 vb_din0[15]
port 277 nsew signal output
rlabel metal3 s 0 71544 800 71664 6 vb_din0[16]
port 278 nsew signal output
rlabel metal3 s 0 74128 800 74248 6 vb_din0[17]
port 279 nsew signal output
rlabel metal3 s 0 76712 800 76832 6 vb_din0[18]
port 280 nsew signal output
rlabel metal3 s 0 79432 800 79552 6 vb_din0[19]
port 281 nsew signal output
rlabel metal3 s 0 10072 800 10192 6 vb_din0[1]
port 282 nsew signal output
rlabel metal3 s 0 82016 800 82136 6 vb_din0[20]
port 283 nsew signal output
rlabel metal3 s 0 84736 800 84856 6 vb_din0[21]
port 284 nsew signal output
rlabel metal3 s 0 87320 800 87440 6 vb_din0[22]
port 285 nsew signal output
rlabel metal3 s 0 89904 800 90024 6 vb_din0[23]
port 286 nsew signal output
rlabel metal3 s 0 92624 800 92744 6 vb_din0[24]
port 287 nsew signal output
rlabel metal3 s 0 95208 800 95328 6 vb_din0[25]
port 288 nsew signal output
rlabel metal3 s 0 97928 800 98048 6 vb_din0[26]
port 289 nsew signal output
rlabel metal3 s 0 100512 800 100632 6 vb_din0[27]
port 290 nsew signal output
rlabel metal3 s 0 103096 800 103216 6 vb_din0[28]
port 291 nsew signal output
rlabel metal3 s 0 105816 800 105936 6 vb_din0[29]
port 292 nsew signal output
rlabel metal3 s 0 15240 800 15360 6 vb_din0[2]
port 293 nsew signal output
rlabel metal3 s 0 108400 800 108520 6 vb_din0[30]
port 294 nsew signal output
rlabel metal3 s 0 110984 800 111104 6 vb_din0[31]
port 295 nsew signal output
rlabel metal3 s 0 20544 800 20664 6 vb_din0[3]
port 296 nsew signal output
rlabel metal3 s 0 25848 800 25968 6 vb_din0[4]
port 297 nsew signal output
rlabel metal3 s 0 30200 800 30320 6 vb_din0[5]
port 298 nsew signal output
rlabel metal3 s 0 34552 800 34672 6 vb_din0[6]
port 299 nsew signal output
rlabel metal3 s 0 39040 800 39160 6 vb_din0[7]
port 300 nsew signal output
rlabel metal3 s 0 43392 800 43512 6 vb_din0[8]
port 301 nsew signal output
rlabel metal3 s 0 47744 800 47864 6 vb_din0[9]
port 302 nsew signal output
rlabel metal3 s 0 5584 800 5704 6 vb_dout0[0]
port 303 nsew signal input
rlabel metal3 s 0 53048 800 53168 6 vb_dout0[10]
port 304 nsew signal input
rlabel metal3 s 0 57400 800 57520 6 vb_dout0[11]
port 305 nsew signal input
rlabel metal3 s 0 61888 800 62008 6 vb_dout0[12]
port 306 nsew signal input
rlabel metal3 s 0 64472 800 64592 6 vb_dout0[13]
port 307 nsew signal input
rlabel metal3 s 0 67056 800 67176 6 vb_dout0[14]
port 308 nsew signal input
rlabel metal3 s 0 69776 800 69896 6 vb_dout0[15]
port 309 nsew signal input
rlabel metal3 s 0 72360 800 72480 6 vb_dout0[16]
port 310 nsew signal input
rlabel metal3 s 0 75080 800 75200 6 vb_dout0[17]
port 311 nsew signal input
rlabel metal3 s 0 77664 800 77784 6 vb_dout0[18]
port 312 nsew signal input
rlabel metal3 s 0 80248 800 80368 6 vb_dout0[19]
port 313 nsew signal input
rlabel metal3 s 0 10888 800 11008 6 vb_dout0[1]
port 314 nsew signal input
rlabel metal3 s 0 82968 800 83088 6 vb_dout0[20]
port 315 nsew signal input
rlabel metal3 s 0 85552 800 85672 6 vb_dout0[21]
port 316 nsew signal input
rlabel metal3 s 0 88136 800 88256 6 vb_dout0[22]
port 317 nsew signal input
rlabel metal3 s 0 90856 800 90976 6 vb_dout0[23]
port 318 nsew signal input
rlabel metal3 s 0 93440 800 93560 6 vb_dout0[24]
port 319 nsew signal input
rlabel metal3 s 0 96160 800 96280 6 vb_dout0[25]
port 320 nsew signal input
rlabel metal3 s 0 98744 800 98864 6 vb_dout0[26]
port 321 nsew signal input
rlabel metal3 s 0 101328 800 101448 6 vb_dout0[27]
port 322 nsew signal input
rlabel metal3 s 0 104048 800 104168 6 vb_dout0[28]
port 323 nsew signal input
rlabel metal3 s 0 106632 800 106752 6 vb_dout0[29]
port 324 nsew signal input
rlabel metal3 s 0 16192 800 16312 6 vb_dout0[2]
port 325 nsew signal input
rlabel metal3 s 0 109216 800 109336 6 vb_dout0[30]
port 326 nsew signal input
rlabel metal3 s 0 111936 800 112056 6 vb_dout0[31]
port 327 nsew signal input
rlabel metal3 s 0 21496 800 21616 6 vb_dout0[3]
port 328 nsew signal input
rlabel metal3 s 0 26664 800 26784 6 vb_dout0[4]
port 329 nsew signal input
rlabel metal3 s 0 31152 800 31272 6 vb_dout0[5]
port 330 nsew signal input
rlabel metal3 s 0 35504 800 35624 6 vb_dout0[6]
port 331 nsew signal input
rlabel metal3 s 0 39856 800 39976 6 vb_dout0[7]
port 332 nsew signal input
rlabel metal3 s 0 44208 800 44328 6 vb_dout0[8]
port 333 nsew signal input
rlabel metal3 s 0 48696 800 48816 6 vb_dout0[9]
port 334 nsew signal input
rlabel metal3 s 0 6536 800 6656 6 vb_dout1[0]
port 335 nsew signal input
rlabel metal3 s 0 54000 800 54120 6 vb_dout1[10]
port 336 nsew signal input
rlabel metal3 s 0 58352 800 58472 6 vb_dout1[11]
port 337 nsew signal input
rlabel metal3 s 0 62704 800 62824 6 vb_dout1[12]
port 338 nsew signal input
rlabel metal3 s 0 65424 800 65544 6 vb_dout1[13]
port 339 nsew signal input
rlabel metal3 s 0 68008 800 68128 6 vb_dout1[14]
port 340 nsew signal input
rlabel metal3 s 0 70592 800 70712 6 vb_dout1[15]
port 341 nsew signal input
rlabel metal3 s 0 73312 800 73432 6 vb_dout1[16]
port 342 nsew signal input
rlabel metal3 s 0 75896 800 76016 6 vb_dout1[17]
port 343 nsew signal input
rlabel metal3 s 0 78480 800 78600 6 vb_dout1[18]
port 344 nsew signal input
rlabel metal3 s 0 81200 800 81320 6 vb_dout1[19]
port 345 nsew signal input
rlabel metal3 s 0 11704 800 11824 6 vb_dout1[1]
port 346 nsew signal input
rlabel metal3 s 0 83784 800 83904 6 vb_dout1[20]
port 347 nsew signal input
rlabel metal3 s 0 86504 800 86624 6 vb_dout1[21]
port 348 nsew signal input
rlabel metal3 s 0 89088 800 89208 6 vb_dout1[22]
port 349 nsew signal input
rlabel metal3 s 0 91672 800 91792 6 vb_dout1[23]
port 350 nsew signal input
rlabel metal3 s 0 94392 800 94512 6 vb_dout1[24]
port 351 nsew signal input
rlabel metal3 s 0 96976 800 97096 6 vb_dout1[25]
port 352 nsew signal input
rlabel metal3 s 0 99560 800 99680 6 vb_dout1[26]
port 353 nsew signal input
rlabel metal3 s 0 102280 800 102400 6 vb_dout1[27]
port 354 nsew signal input
rlabel metal3 s 0 104864 800 104984 6 vb_dout1[28]
port 355 nsew signal input
rlabel metal3 s 0 107584 800 107704 6 vb_dout1[29]
port 356 nsew signal input
rlabel metal3 s 0 17008 800 17128 6 vb_dout1[2]
port 357 nsew signal input
rlabel metal3 s 0 110168 800 110288 6 vb_dout1[30]
port 358 nsew signal input
rlabel metal3 s 0 112752 800 112872 6 vb_dout1[31]
port 359 nsew signal input
rlabel metal3 s 0 22312 800 22432 6 vb_dout1[3]
port 360 nsew signal input
rlabel metal3 s 0 27616 800 27736 6 vb_dout1[4]
port 361 nsew signal input
rlabel metal3 s 0 31968 800 32088 6 vb_dout1[5]
port 362 nsew signal input
rlabel metal3 s 0 36320 800 36440 6 vb_dout1[6]
port 363 nsew signal input
rlabel metal3 s 0 40808 800 40928 6 vb_dout1[7]
port 364 nsew signal input
rlabel metal3 s 0 45160 800 45280 6 vb_dout1[8]
port 365 nsew signal input
rlabel metal3 s 0 49512 800 49632 6 vb_dout1[9]
port 366 nsew signal input
rlabel metal3 s 0 2048 800 2168 6 vb_web0
port 367 nsew signal output
rlabel metal3 s 0 7352 800 7472 6 vb_wmask0[0]
port 368 nsew signal output
rlabel metal3 s 0 12656 800 12776 6 vb_wmask0[1]
port 369 nsew signal output
rlabel metal3 s 0 17960 800 18080 6 vb_wmask0[2]
port 370 nsew signal output
rlabel metal3 s 0 23128 800 23248 6 vb_wmask0[3]
port 371 nsew signal output
rlabel metal4 s 4208 2128 4528 257360 6 vccd1
port 372 nsew power input
rlabel metal4 s 34928 2128 35248 257360 6 vccd1
port 372 nsew power input
rlabel metal4 s 65648 2128 65968 257360 6 vccd1
port 372 nsew power input
rlabel metal4 s 96368 2128 96688 257360 6 vccd1
port 372 nsew power input
rlabel metal4 s 127088 2128 127408 257360 6 vccd1
port 372 nsew power input
rlabel metal4 s 157808 2128 158128 257360 6 vccd1
port 372 nsew power input
rlabel metal4 s 188528 2128 188848 257360 6 vccd1
port 372 nsew power input
rlabel metal4 s 219248 2128 219568 257360 6 vccd1
port 372 nsew power input
rlabel metal4 s 249968 2128 250288 257360 6 vccd1
port 372 nsew power input
rlabel metal4 s 19568 2128 19888 257360 6 vssd1
port 373 nsew ground input
rlabel metal4 s 50288 2128 50608 257360 6 vssd1
port 373 nsew ground input
rlabel metal4 s 81008 2128 81328 257360 6 vssd1
port 373 nsew ground input
rlabel metal4 s 111728 2128 112048 257360 6 vssd1
port 373 nsew ground input
rlabel metal4 s 142448 2128 142768 257360 6 vssd1
port 373 nsew ground input
rlabel metal4 s 173168 2128 173488 257360 6 vssd1
port 373 nsew ground input
rlabel metal4 s 203888 2128 204208 257360 6 vssd1
port 373 nsew ground input
rlabel metal4 s 234608 2128 234928 257360 6 vssd1
port 373 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 260000 260000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 70259250
string GDS_FILE /home/kasirga/c0_hayyan/GL_GECTI/caravel_user_project/openlane/c0_system/runs/c0_system/results/finishing/c0_system.magic.gds
string GDS_START 1649888
<< end >>


magic
tech sky130A
magscale 1 2
timestamp 1647619795
<< metal1 >>
rect 201494 702992 201500 703044
rect 201552 703032 201558 703044
rect 202782 703032 202788 703044
rect 201552 703004 202788 703032
rect 201552 702992 201558 703004
rect 202782 702992 202788 703004
rect 202840 702992 202846 703044
rect 413646 700476 413652 700528
rect 413704 700516 413710 700528
rect 420914 700516 420920 700528
rect 413704 700488 420920 700516
rect 413704 700476 413710 700488
rect 420914 700476 420920 700488
rect 420972 700476 420978 700528
rect 154114 700340 154120 700392
rect 154172 700380 154178 700392
rect 189718 700380 189724 700392
rect 154172 700352 189724 700380
rect 154172 700340 154178 700352
rect 189718 700340 189724 700352
rect 189776 700340 189782 700392
rect 278774 700340 278780 700392
rect 278832 700380 278838 700392
rect 348786 700380 348792 700392
rect 278832 700352 348792 700380
rect 278832 700340 278838 700352
rect 348786 700340 348792 700352
rect 348844 700340 348850 700392
rect 72970 700272 72976 700324
rect 73028 700312 73034 700324
rect 239398 700312 239404 700324
rect 73028 700284 239404 700312
rect 73028 700272 73034 700284
rect 239398 700272 239404 700284
rect 239456 700272 239462 700324
rect 262214 700272 262220 700324
rect 262272 700312 262278 700324
rect 332502 700312 332508 700324
rect 262272 700284 332508 700312
rect 262272 700272 262278 700284
rect 332502 700272 332508 700284
rect 332560 700272 332566 700324
rect 527174 700272 527180 700324
rect 527232 700312 527238 700324
rect 538214 700312 538220 700324
rect 527232 700284 538220 700312
rect 527232 700272 527238 700284
rect 538214 700272 538220 700284
rect 538272 700272 538278 700324
rect 397454 699932 397460 699984
rect 397512 699972 397518 699984
rect 399294 699972 399300 699984
rect 397512 699944 399300 699972
rect 397512 699932 397518 699944
rect 399294 699932 399300 699944
rect 399352 699932 399358 699984
rect 266354 697552 266360 697604
rect 266412 697592 266418 697604
rect 267642 697592 267648 697604
rect 266412 697564 267648 697592
rect 266412 697552 266418 697564
rect 267642 697552 267648 697564
rect 267700 697552 267706 697604
rect 399294 695444 399300 695496
rect 399352 695484 399358 695496
rect 400950 695484 400956 695496
rect 399352 695456 400956 695484
rect 399352 695444 399358 695456
rect 400950 695444 400956 695456
rect 401008 695444 401014 695496
rect 477494 694764 477500 694816
rect 477552 694804 477558 694816
rect 480254 694804 480260 694816
rect 477552 694776 480260 694804
rect 477552 694764 477558 694776
rect 480254 694764 480260 694776
rect 480312 694764 480318 694816
rect 420914 694152 420920 694204
rect 420972 694192 420978 694204
rect 424318 694192 424324 694204
rect 420972 694164 424324 694192
rect 420972 694152 420978 694164
rect 424318 694152 424324 694164
rect 424376 694152 424382 694204
rect 259454 694084 259460 694136
rect 259512 694124 259518 694136
rect 262122 694124 262128 694136
rect 259512 694096 262128 694124
rect 259512 694084 259518 694096
rect 262122 694084 262128 694096
rect 262180 694084 262186 694136
rect 276750 692792 276756 692844
rect 276808 692832 276814 692844
rect 278682 692832 278688 692844
rect 276808 692804 278688 692832
rect 276808 692792 276814 692804
rect 278682 692792 278688 692804
rect 278740 692792 278746 692844
rect 400950 691092 400956 691144
rect 401008 691132 401014 691144
rect 401962 691132 401968 691144
rect 401008 691104 401968 691132
rect 401008 691092 401014 691104
rect 401962 691092 401968 691104
rect 402020 691092 402026 691144
rect 462314 690684 462320 690736
rect 462372 690724 462378 690736
rect 465166 690724 465172 690736
rect 462372 690696 465172 690724
rect 462372 690684 462378 690696
rect 465166 690684 465172 690696
rect 465224 690684 465230 690736
rect 465166 688168 465172 688220
rect 465224 688208 465230 688220
rect 471238 688208 471244 688220
rect 465224 688180 471244 688208
rect 465224 688168 465230 688180
rect 471238 688168 471244 688180
rect 471296 688168 471302 688220
rect 480254 687896 480260 687948
rect 480312 687936 480318 687948
rect 490558 687936 490564 687948
rect 480312 687908 490564 687936
rect 480312 687896 480318 687908
rect 490558 687896 490564 687908
rect 490616 687896 490622 687948
rect 275278 687488 275284 687540
rect 275336 687528 275342 687540
rect 276750 687528 276756 687540
rect 275336 687500 276756 687528
rect 275336 687488 275342 687500
rect 276750 687488 276756 687500
rect 276808 687488 276814 687540
rect 424318 685108 424324 685160
rect 424376 685148 424382 685160
rect 447778 685148 447784 685160
rect 424376 685120 447784 685148
rect 424376 685108 424382 685120
rect 447778 685108 447784 685120
rect 447836 685108 447842 685160
rect 401962 684496 401968 684548
rect 402020 684536 402026 684548
rect 402020 684508 402974 684536
rect 402020 684496 402026 684508
rect 402946 684468 402974 684508
rect 404998 684468 405004 684480
rect 402946 684440 405004 684468
rect 404998 684428 405004 684440
rect 405056 684428 405062 684480
rect 253198 683136 253204 683188
rect 253256 683176 253262 683188
rect 259362 683176 259368 683188
rect 253256 683148 259368 683176
rect 253256 683136 253262 683148
rect 259362 683136 259368 683148
rect 259420 683136 259426 683188
rect 471238 681368 471244 681420
rect 471296 681408 471302 681420
rect 474642 681408 474648 681420
rect 471296 681380 474648 681408
rect 471296 681368 471302 681380
rect 474642 681368 474648 681380
rect 474700 681368 474706 681420
rect 474642 677492 474648 677544
rect 474700 677532 474706 677544
rect 478138 677532 478144 677544
rect 474700 677504 478144 677532
rect 474700 677492 474706 677504
rect 478138 677492 478144 677504
rect 478196 677492 478202 677544
rect 478138 672732 478144 672784
rect 478196 672772 478202 672784
rect 483658 672772 483664 672784
rect 478196 672744 483664 672772
rect 478196 672732 478202 672744
rect 483658 672732 483664 672744
rect 483716 672732 483722 672784
rect 490558 665116 490564 665168
rect 490616 665156 490622 665168
rect 493318 665156 493324 665168
rect 490616 665128 493324 665156
rect 490616 665116 490622 665128
rect 493318 665116 493324 665128
rect 493376 665116 493382 665168
rect 447778 664436 447784 664488
rect 447836 664476 447842 664488
rect 460198 664476 460204 664488
rect 447836 664448 460204 664476
rect 447836 664436 447842 664448
rect 460198 664436 460204 664448
rect 460256 664436 460262 664488
rect 483658 664436 483664 664488
rect 483716 664476 483722 664488
rect 497458 664476 497464 664488
rect 483716 664448 497464 664476
rect 483716 664436 483722 664448
rect 497458 664436 497464 664448
rect 497516 664436 497522 664488
rect 3510 656888 3516 656940
rect 3568 656928 3574 656940
rect 239582 656928 239588 656940
rect 3568 656900 239588 656928
rect 3568 656888 3574 656900
rect 239582 656888 239588 656900
rect 239640 656888 239646 656940
rect 460198 656276 460204 656328
rect 460256 656316 460262 656328
rect 462314 656316 462320 656328
rect 460256 656288 462320 656316
rect 460256 656276 460262 656288
rect 462314 656276 462320 656288
rect 462372 656276 462378 656328
rect 273898 655460 273904 655512
rect 273956 655500 273962 655512
rect 275278 655500 275284 655512
rect 273956 655472 275284 655500
rect 273956 655460 273962 655472
rect 275278 655460 275284 655472
rect 275336 655460 275342 655512
rect 497458 654780 497464 654832
rect 497516 654820 497522 654832
rect 508498 654820 508504 654832
rect 497516 654792 508504 654820
rect 497516 654780 497522 654792
rect 508498 654780 508504 654792
rect 508556 654780 508562 654832
rect 462314 653148 462320 653200
rect 462372 653188 462378 653200
rect 465442 653188 465448 653200
rect 462372 653160 465448 653188
rect 462372 653148 462378 653160
rect 465442 653148 465448 653160
rect 465500 653148 465506 653200
rect 465442 650632 465448 650684
rect 465500 650672 465506 650684
rect 480898 650672 480904 650684
rect 465500 650644 480904 650672
rect 465500 650632 465506 650644
rect 480898 650632 480904 650644
rect 480956 650632 480962 650684
rect 480898 641044 480904 641096
rect 480956 641084 480962 641096
rect 494698 641084 494704 641096
rect 480956 641056 494704 641084
rect 480956 641044 480962 641056
rect 494698 641044 494704 641056
rect 494756 641044 494762 641096
rect 493318 640976 493324 641028
rect 493376 641016 493382 641028
rect 507118 641016 507124 641028
rect 493376 640988 507124 641016
rect 493376 640976 493382 640988
rect 507118 640976 507124 640988
rect 507176 640976 507182 641028
rect 272518 638188 272524 638240
rect 272576 638228 272582 638240
rect 273898 638228 273904 638240
rect 272576 638200 273904 638228
rect 272576 638188 272582 638200
rect 273898 638188 273904 638200
rect 273956 638188 273962 638240
rect 494698 636828 494704 636880
rect 494756 636868 494762 636880
rect 505738 636868 505744 636880
rect 494756 636840 505744 636868
rect 494756 636828 494762 636840
rect 505738 636828 505744 636840
rect 505796 636828 505802 636880
rect 508498 633700 508504 633752
rect 508556 633740 508562 633752
rect 511258 633740 511264 633752
rect 508556 633712 511264 633740
rect 508556 633700 508562 633712
rect 511258 633700 511264 633712
rect 511316 633700 511322 633752
rect 251818 627852 251824 627904
rect 251876 627892 251882 627904
rect 253198 627892 253204 627904
rect 251876 627864 253204 627892
rect 251876 627852 251882 627864
rect 253198 627852 253204 627864
rect 253256 627852 253262 627904
rect 404998 626492 405004 626544
rect 405056 626532 405062 626544
rect 407758 626532 407764 626544
rect 405056 626504 407764 626532
rect 405056 626492 405062 626504
rect 407758 626492 407764 626504
rect 407816 626492 407822 626544
rect 511258 624384 511264 624436
rect 511316 624424 511322 624436
rect 521654 624424 521660 624436
rect 511316 624396 521660 624424
rect 511316 624384 511322 624396
rect 521654 624384 521660 624396
rect 521712 624384 521718 624436
rect 269758 623772 269764 623824
rect 269816 623812 269822 623824
rect 272518 623812 272524 623824
rect 269816 623784 272524 623812
rect 269816 623772 269822 623784
rect 272518 623772 272524 623784
rect 272576 623772 272582 623824
rect 505738 623024 505744 623076
rect 505796 623064 505802 623076
rect 522298 623064 522304 623076
rect 505796 623036 522304 623064
rect 505796 623024 505802 623036
rect 522298 623024 522304 623036
rect 522356 623024 522362 623076
rect 521654 616768 521660 616820
rect 521712 616808 521718 616820
rect 525150 616808 525156 616820
rect 521712 616780 525156 616808
rect 521712 616768 521718 616780
rect 525150 616768 525156 616780
rect 525208 616768 525214 616820
rect 522298 614184 522304 614236
rect 522356 614224 522362 614236
rect 525058 614224 525064 614236
rect 522356 614196 525064 614224
rect 522356 614184 522362 614196
rect 525058 614184 525064 614196
rect 525116 614184 525122 614236
rect 407758 613028 407764 613080
rect 407816 613068 407822 613080
rect 409230 613068 409236 613080
rect 407816 613040 409236 613068
rect 407816 613028 407822 613040
rect 409230 613028 409236 613040
rect 409288 613028 409294 613080
rect 409230 609900 409236 609952
rect 409288 609940 409294 609952
rect 410518 609940 410524 609952
rect 409288 609912 410524 609940
rect 409288 609900 409294 609912
rect 410518 609900 410524 609912
rect 410576 609900 410582 609952
rect 507118 607860 507124 607912
rect 507176 607900 507182 607912
rect 518894 607900 518900 607912
rect 507176 607872 518900 607900
rect 507176 607860 507182 607872
rect 518894 607860 518900 607872
rect 518952 607860 518958 607912
rect 525150 607112 525156 607164
rect 525208 607152 525214 607164
rect 527634 607152 527640 607164
rect 525208 607124 527640 607152
rect 525208 607112 525214 607124
rect 527634 607112 527640 607124
rect 527692 607112 527698 607164
rect 268746 604460 268752 604512
rect 268804 604500 268810 604512
rect 269758 604500 269764 604512
rect 268804 604472 269764 604500
rect 268804 604460 268810 604472
rect 269758 604460 269764 604472
rect 269816 604460 269822 604512
rect 527634 603712 527640 603764
rect 527692 603752 527698 603764
rect 533338 603752 533344 603764
rect 527692 603724 533344 603752
rect 527692 603712 527698 603724
rect 533338 603712 533344 603724
rect 533396 603712 533402 603764
rect 518894 603100 518900 603152
rect 518952 603140 518958 603152
rect 522850 603140 522856 603152
rect 518952 603112 522856 603140
rect 518952 603100 518958 603112
rect 522850 603100 522856 603112
rect 522908 603100 522914 603152
rect 266998 602352 267004 602404
rect 267056 602392 267062 602404
rect 268746 602392 268752 602404
rect 267056 602364 268752 602392
rect 267056 602352 267062 602364
rect 268746 602352 268752 602364
rect 268804 602352 268810 602404
rect 250438 600448 250444 600500
rect 250496 600488 250502 600500
rect 251818 600488 251824 600500
rect 250496 600460 251824 600488
rect 250496 600448 250502 600460
rect 251818 600448 251824 600460
rect 251876 600448 251882 600500
rect 410518 600244 410524 600296
rect 410576 600284 410582 600296
rect 411898 600284 411904 600296
rect 410576 600256 411904 600284
rect 410576 600244 410582 600256
rect 411898 600244 411904 600256
rect 411956 600244 411962 600296
rect 411898 595076 411904 595128
rect 411956 595116 411962 595128
rect 414658 595116 414664 595128
rect 411956 595088 414664 595116
rect 411956 595076 411962 595088
rect 414658 595076 414664 595088
rect 414716 595076 414722 595128
rect 533338 591948 533344 592000
rect 533396 591988 533402 592000
rect 538306 591988 538312 592000
rect 533396 591960 538312 591988
rect 533396 591948 533402 591960
rect 538306 591948 538312 591960
rect 538364 591948 538370 592000
rect 282178 588412 282184 588464
rect 282236 588452 282242 588464
rect 282914 588452 282920 588464
rect 282236 588424 282920 588452
rect 282236 588412 282242 588424
rect 282914 588412 282920 588424
rect 282972 588412 282978 588464
rect 264974 579640 264980 579692
rect 265032 579680 265038 579692
rect 266998 579680 267004 579692
rect 265032 579652 267004 579680
rect 265032 579640 265038 579652
rect 266998 579640 267004 579652
rect 267056 579640 267062 579692
rect 262858 578144 262864 578196
rect 262916 578184 262922 578196
rect 264974 578184 264980 578196
rect 262916 578156 264980 578184
rect 262916 578144 262922 578156
rect 264974 578144 264980 578156
rect 265032 578144 265038 578196
rect 577498 577192 577504 577244
rect 577556 577232 577562 577244
rect 579614 577232 579620 577244
rect 577556 577204 579620 577232
rect 577556 577192 577562 577204
rect 579614 577192 579620 577204
rect 579672 577192 579678 577244
rect 280798 575492 280804 575544
rect 280856 575532 280862 575544
rect 282178 575532 282184 575544
rect 280856 575504 282184 575532
rect 280856 575492 280862 575504
rect 282178 575492 282184 575504
rect 282236 575492 282242 575544
rect 247678 573792 247684 573844
rect 247736 573832 247742 573844
rect 250438 573832 250444 573844
rect 247736 573804 250444 573832
rect 247736 573792 247742 573804
rect 250438 573792 250444 573804
rect 250496 573792 250502 573844
rect 3050 565836 3056 565888
rect 3108 565876 3114 565888
rect 191098 565876 191104 565888
rect 3108 565848 191104 565876
rect 3108 565836 3114 565848
rect 191098 565836 191104 565848
rect 191156 565836 191162 565888
rect 525058 562300 525064 562352
rect 525116 562340 525122 562352
rect 533338 562340 533344 562352
rect 525116 562312 533344 562340
rect 525116 562300 525122 562312
rect 533338 562300 533344 562312
rect 533396 562300 533402 562352
rect 280798 561728 280804 561740
rect 278792 561700 280804 561728
rect 278038 561620 278044 561672
rect 278096 561660 278102 561672
rect 278792 561660 278820 561700
rect 280798 561688 280804 561700
rect 280856 561688 280862 561740
rect 278096 561632 278820 561660
rect 278096 561620 278102 561632
rect 414658 558832 414664 558884
rect 414716 558872 414722 558884
rect 416038 558872 416044 558884
rect 414716 558844 416044 558872
rect 414716 558832 414722 558844
rect 416038 558832 416044 558844
rect 416096 558832 416102 558884
rect 3602 553392 3608 553444
rect 3660 553432 3666 553444
rect 239766 553432 239772 553444
rect 3660 553404 239772 553432
rect 3660 553392 3666 553404
rect 239766 553392 239772 553404
rect 239824 553392 239830 553444
rect 261202 550740 261208 550792
rect 261260 550780 261266 550792
rect 262858 550780 262864 550792
rect 261260 550752 262864 550780
rect 261260 550740 261266 550752
rect 262858 550740 262864 550752
rect 262916 550740 262922 550792
rect 259454 548496 259460 548548
rect 259512 548536 259518 548548
rect 261202 548536 261208 548548
rect 259512 548508 261208 548536
rect 259512 548496 259518 548508
rect 261202 548496 261208 548508
rect 261260 548496 261266 548548
rect 533338 543804 533344 543856
rect 533396 543844 533402 543856
rect 535730 543844 535736 543856
rect 533396 543816 535736 543844
rect 533396 543804 533402 543816
rect 535730 543804 535736 543816
rect 535788 543804 535794 543856
rect 535730 542308 535736 542360
rect 535788 542348 535794 542360
rect 538030 542348 538036 542360
rect 535788 542320 538036 542348
rect 535788 542308 535794 542320
rect 538030 542308 538036 542320
rect 538088 542308 538094 542360
rect 257338 539588 257344 539640
rect 257396 539628 257402 539640
rect 259362 539628 259368 539640
rect 257396 539600 259368 539628
rect 257396 539588 257402 539600
rect 259362 539588 259368 539600
rect 259420 539588 259426 539640
rect 245010 532448 245016 532500
rect 245068 532488 245074 532500
rect 247678 532488 247684 532500
rect 245068 532460 247684 532488
rect 245068 532448 245074 532460
rect 247678 532448 247684 532460
rect 247736 532448 247742 532500
rect 416038 529864 416044 529916
rect 416096 529904 416102 529916
rect 417510 529904 417516 529916
rect 416096 529876 417516 529904
rect 416096 529864 416102 529876
rect 417510 529864 417516 529876
rect 417568 529864 417574 529916
rect 417510 526260 417516 526312
rect 417568 526300 417574 526312
rect 418890 526300 418896 526312
rect 417568 526272 418896 526300
rect 417568 526260 417574 526272
rect 418890 526260 418896 526272
rect 418948 526260 418954 526312
rect 254578 524424 254584 524476
rect 254636 524464 254642 524476
rect 257338 524464 257344 524476
rect 254636 524436 257344 524464
rect 254636 524424 254642 524436
rect 257338 524424 257344 524436
rect 257396 524424 257402 524476
rect 577590 524424 577596 524476
rect 577648 524464 577654 524476
rect 579614 524464 579620 524476
rect 577648 524436 579620 524464
rect 577648 524424 577654 524436
rect 579614 524424 579620 524436
rect 579672 524424 579678 524476
rect 244918 523676 244924 523728
rect 244976 523716 244982 523728
rect 278038 523716 278044 523728
rect 244976 523688 278044 523716
rect 244976 523676 244982 523688
rect 278038 523676 278044 523688
rect 278096 523676 278102 523728
rect 418890 521568 418896 521620
rect 418948 521608 418954 521620
rect 420178 521608 420184 521620
rect 418948 521580 420184 521608
rect 418948 521568 418954 521580
rect 420178 521568 420184 521580
rect 420236 521568 420242 521620
rect 3326 514768 3332 514820
rect 3384 514808 3390 514820
rect 235258 514808 235264 514820
rect 3384 514780 235264 514808
rect 3384 514768 3390 514780
rect 235258 514768 235264 514780
rect 235316 514768 235322 514820
rect 420178 514700 420184 514752
rect 420236 514740 420242 514752
rect 422938 514740 422944 514752
rect 420236 514712 422944 514740
rect 420236 514700 420242 514712
rect 422938 514700 422944 514712
rect 422996 514700 423002 514752
rect 243630 506472 243636 506524
rect 243688 506512 243694 506524
rect 245010 506512 245016 506524
rect 243688 506484 245016 506512
rect 243688 506472 243694 506484
rect 245010 506472 245016 506484
rect 245068 506472 245074 506524
rect 422938 505724 422944 505776
rect 422996 505764 423002 505776
rect 424318 505764 424324 505776
rect 422996 505736 424324 505764
rect 422996 505724 423002 505736
rect 424318 505724 424324 505736
rect 424376 505724 424382 505776
rect 251634 505112 251640 505164
rect 251692 505152 251698 505164
rect 254578 505152 254584 505164
rect 251692 505124 254584 505152
rect 251692 505112 251698 505124
rect 254578 505112 254584 505124
rect 254636 505112 254642 505164
rect 242158 504160 242164 504212
rect 242216 504200 242222 504212
rect 243630 504200 243636 504212
rect 242216 504172 243636 504200
rect 242216 504160 242222 504172
rect 243630 504160 243636 504172
rect 243688 504160 243694 504212
rect 249794 501984 249800 502036
rect 249852 502024 249858 502036
rect 251634 502024 251640 502036
rect 249852 501996 251640 502024
rect 249852 501984 249858 501996
rect 251634 501984 251640 501996
rect 251692 501984 251698 502036
rect 3326 500964 3332 501016
rect 3384 501004 3390 501016
rect 239490 501004 239496 501016
rect 3384 500976 239496 501004
rect 3384 500964 3390 500976
rect 239490 500964 239496 500976
rect 239548 500964 239554 501016
rect 247678 496952 247684 497004
rect 247736 496992 247742 497004
rect 249794 496992 249800 497004
rect 247736 496964 249800 496992
rect 247736 496952 247742 496964
rect 249794 496952 249800 496964
rect 249852 496952 249858 497004
rect 242250 496816 242256 496868
rect 242308 496856 242314 496868
rect 244918 496856 244924 496868
rect 242308 496828 244924 496856
rect 242308 496816 242314 496828
rect 244918 496816 244924 496828
rect 244976 496816 244982 496868
rect 242802 485800 242808 485852
rect 242860 485840 242866 485852
rect 247678 485840 247684 485852
rect 242860 485812 247684 485840
rect 242860 485800 242866 485812
rect 247678 485800 247684 485812
rect 247736 485800 247742 485852
rect 240318 484032 240324 484084
rect 240376 484072 240382 484084
rect 242250 484072 242256 484084
rect 240376 484044 242256 484072
rect 240376 484032 240382 484044
rect 242250 484032 242256 484044
rect 242308 484032 242314 484084
rect 240778 483760 240784 483812
rect 240836 483800 240842 483812
rect 242802 483800 242808 483812
rect 240836 483772 242808 483800
rect 240836 483760 240842 483772
rect 242802 483760 242808 483772
rect 242860 483760 242866 483812
rect 239858 482672 239864 482724
rect 239916 482712 239922 482724
rect 242158 482712 242164 482724
rect 239916 482684 242164 482712
rect 239916 482672 239922 482684
rect 242158 482672 242164 482684
rect 242216 482672 242222 482724
rect 239674 480904 239680 480956
rect 239732 480944 239738 480956
rect 266354 480944 266360 480956
rect 239732 480916 266360 480944
rect 239732 480904 239738 480916
rect 266354 480904 266360 480916
rect 266412 480904 266418 480956
rect 424318 480904 424324 480956
rect 424376 480944 424382 480956
rect 437382 480944 437388 480956
rect 424376 480916 437388 480944
rect 424376 480904 424382 480916
rect 437382 480904 437388 480916
rect 437440 480904 437446 480956
rect 239214 479544 239220 479596
rect 239272 479584 239278 479596
rect 240778 479584 240784 479596
rect 239272 479556 240784 479584
rect 239272 479544 239278 479556
rect 240778 479544 240784 479556
rect 240836 479544 240842 479596
rect 437382 479544 437388 479596
rect 437440 479544 437446 479596
rect 437400 479516 437428 479544
rect 538398 479516 538404 479528
rect 437400 479488 538404 479516
rect 538398 479476 538404 479488
rect 538456 479476 538462 479528
rect 157242 478864 157248 478916
rect 157300 478904 157306 478916
rect 237374 478904 237380 478916
rect 157300 478876 237380 478904
rect 157300 478864 157306 478876
rect 237374 478864 237380 478876
rect 237432 478864 237438 478916
rect 239306 478864 239312 478916
rect 239364 478904 239370 478916
rect 240318 478904 240324 478916
rect 239364 478876 240324 478904
rect 239364 478864 239370 478876
rect 240318 478864 240324 478876
rect 240376 478864 240382 478916
rect 235534 477504 235540 477556
rect 235592 477544 235598 477556
rect 237374 477544 237380 477556
rect 235592 477516 237380 477544
rect 235592 477504 235598 477516
rect 237374 477504 237380 477516
rect 237432 477504 237438 477556
rect 235626 476076 235632 476128
rect 235684 476116 235690 476128
rect 237374 476116 237380 476128
rect 235684 476088 237380 476116
rect 235684 476076 235690 476088
rect 237374 476076 237380 476088
rect 237432 476076 237438 476128
rect 154482 473356 154488 473408
rect 154540 473396 154546 473408
rect 237374 473396 237380 473408
rect 154540 473368 237380 473396
rect 154540 473356 154546 473368
rect 237374 473356 237380 473368
rect 237432 473356 237438 473408
rect 235718 472064 235724 472116
rect 235776 472104 235782 472116
rect 237466 472104 237472 472116
rect 235776 472076 237472 472104
rect 235776 472064 235782 472076
rect 237466 472064 237472 472076
rect 237524 472064 237530 472116
rect 235810 471996 235816 472048
rect 235868 472036 235874 472048
rect 237374 472036 237380 472048
rect 235868 472008 237380 472036
rect 235868 471996 235874 472008
rect 237374 471996 237380 472008
rect 237432 471996 237438 472048
rect 151354 469208 151360 469260
rect 151412 469248 151418 469260
rect 237374 469248 237380 469260
rect 151412 469220 237380 469248
rect 151412 469208 151418 469220
rect 237374 469208 237380 469220
rect 237432 469208 237438 469260
rect 235902 467848 235908 467900
rect 235960 467888 235966 467900
rect 237374 467888 237380 467900
rect 235960 467860 237380 467888
rect 235960 467848 235966 467860
rect 237374 467848 237380 467860
rect 237432 467848 237438 467900
rect 235166 466420 235172 466472
rect 235224 466460 235230 466472
rect 237374 466460 237380 466472
rect 235224 466432 237380 466460
rect 235224 466420 235230 466432
rect 237374 466420 237380 466432
rect 237432 466420 237438 466472
rect 169754 465944 169760 465996
rect 169812 465984 169818 465996
rect 192478 465984 192484 465996
rect 169812 465956 192484 465984
rect 169812 465944 169818 465956
rect 192478 465944 192484 465956
rect 192536 465944 192542 465996
rect 168466 465876 168472 465928
rect 168524 465916 168530 465928
rect 192570 465916 192576 465928
rect 168524 465888 192576 465916
rect 168524 465876 168530 465888
rect 192570 465876 192576 465888
rect 192628 465876 192634 465928
rect 146018 465808 146024 465860
rect 146076 465848 146082 465860
rect 186682 465848 186688 465860
rect 146076 465820 186688 465848
rect 146076 465808 146082 465820
rect 186682 465808 186688 465820
rect 186740 465808 186746 465860
rect 141050 465740 141056 465792
rect 141108 465780 141114 465792
rect 187234 465780 187240 465792
rect 141108 465752 187240 465780
rect 141108 465740 141114 465752
rect 187234 465740 187240 465752
rect 187292 465740 187298 465792
rect 136082 465672 136088 465724
rect 136140 465712 136146 465724
rect 187142 465712 187148 465724
rect 136140 465684 187148 465712
rect 136140 465672 136146 465684
rect 187142 465672 187148 465684
rect 187200 465672 187206 465724
rect 128722 465604 128728 465656
rect 128780 465644 128786 465656
rect 187050 465644 187056 465656
rect 128780 465616 187056 465644
rect 128780 465604 128786 465616
rect 187050 465604 187056 465616
rect 187108 465604 187114 465656
rect 111058 465536 111064 465588
rect 111116 465576 111122 465588
rect 186958 465576 186964 465588
rect 111116 465548 186964 465576
rect 111116 465536 111122 465548
rect 186958 465536 186964 465548
rect 187016 465536 187022 465588
rect 108482 465468 108488 465520
rect 108540 465508 108546 465520
rect 188338 465508 188344 465520
rect 108540 465480 188344 465508
rect 108540 465468 108546 465480
rect 188338 465468 188344 465480
rect 188396 465468 188402 465520
rect 101306 465400 101312 465452
rect 101364 465440 101370 465452
rect 191282 465440 191288 465452
rect 101364 465412 191288 465440
rect 101364 465400 101370 465412
rect 191282 465400 191288 465412
rect 191340 465400 191346 465452
rect 106182 465332 106188 465384
rect 106240 465372 106246 465384
rect 198182 465372 198188 465384
rect 106240 465344 198188 465372
rect 106240 465332 106246 465344
rect 198182 465332 198188 465344
rect 198240 465332 198246 465384
rect 103698 465264 103704 465316
rect 103756 465304 103762 465316
rect 198090 465304 198096 465316
rect 103756 465276 198096 465304
rect 103756 465264 103762 465276
rect 198090 465264 198096 465276
rect 198148 465264 198154 465316
rect 96154 465196 96160 465248
rect 96212 465236 96218 465248
rect 191190 465236 191196 465248
rect 96212 465208 191196 465236
rect 96212 465196 96218 465208
rect 191190 465196 191196 465208
rect 191248 465196 191254 465248
rect 93670 465128 93676 465180
rect 93728 465168 93734 465180
rect 197998 465168 198004 465180
rect 93728 465140 198004 465168
rect 93728 465128 93734 465140
rect 197998 465128 198004 465140
rect 198056 465128 198062 465180
rect 91186 465060 91192 465112
rect 91244 465100 91250 465112
rect 235442 465100 235448 465112
rect 91244 465072 235448 465100
rect 91244 465060 91250 465072
rect 235442 465060 235448 465072
rect 235500 465060 235506 465112
rect 148502 464992 148508 465044
rect 148560 465032 148566 465044
rect 237374 465032 237380 465044
rect 148560 465004 237380 465032
rect 148560 464992 148566 465004
rect 237374 464992 237380 465004
rect 237432 464992 237438 465044
rect 120994 464924 121000 464976
rect 121052 464964 121058 464976
rect 189902 464964 189908 464976
rect 121052 464936 189908 464964
rect 121052 464924 121058 464936
rect 189902 464924 189908 464936
rect 189960 464924 189966 464976
rect 143626 464856 143632 464908
rect 143684 464896 143690 464908
rect 238018 464896 238024 464908
rect 143684 464868 238024 464896
rect 143684 464856 143690 464868
rect 238018 464856 238024 464868
rect 238076 464856 238082 464908
rect 98546 464788 98552 464840
rect 98604 464828 98610 464840
rect 199378 464828 199384 464840
rect 98604 464800 199384 464828
rect 98604 464788 98610 464800
rect 199378 464788 199384 464800
rect 199436 464788 199442 464840
rect 133506 464720 133512 464772
rect 133564 464760 133570 464772
rect 237926 464760 237932 464772
rect 133564 464732 237932 464760
rect 133564 464720 133570 464732
rect 237926 464720 237932 464732
rect 237984 464720 237990 464772
rect 131114 464652 131120 464704
rect 131172 464692 131178 464704
rect 238662 464692 238668 464704
rect 131172 464664 238668 464692
rect 131172 464652 131178 464664
rect 238662 464652 238668 464664
rect 238720 464652 238726 464704
rect 88518 464584 88524 464636
rect 88576 464624 88582 464636
rect 196618 464624 196624 464636
rect 88576 464596 196624 464624
rect 88576 464584 88582 464596
rect 196618 464584 196624 464596
rect 196676 464584 196682 464636
rect 83458 464516 83464 464568
rect 83516 464556 83522 464568
rect 193858 464556 193864 464568
rect 83516 464528 193864 464556
rect 83516 464516 83522 464528
rect 193858 464516 193864 464528
rect 193916 464516 193922 464568
rect 118602 464448 118608 464500
rect 118660 464488 118666 464500
rect 238386 464488 238392 464500
rect 118660 464460 238392 464488
rect 118660 464448 118666 464460
rect 238386 464448 238392 464460
rect 238444 464448 238450 464500
rect 116118 464380 116124 464432
rect 116176 464420 116182 464432
rect 238202 464420 238208 464432
rect 116176 464392 238208 464420
rect 116176 464380 116182 464392
rect 238202 464380 238208 464392
rect 238260 464380 238266 464432
rect 113634 464312 113640 464364
rect 113692 464352 113698 464364
rect 238110 464352 238116 464364
rect 113692 464324 238116 464352
rect 113692 464312 113698 464324
rect 238110 464312 238116 464324
rect 238168 464312 238174 464364
rect 123570 464244 123576 464296
rect 123628 464284 123634 464296
rect 190086 464284 190092 464296
rect 123628 464256 190092 464284
rect 123628 464244 123634 464256
rect 190086 464244 190092 464256
rect 190144 464244 190150 464296
rect 125962 464176 125968 464228
rect 126020 464216 126026 464228
rect 192662 464216 192668 464228
rect 126020 464188 192668 464216
rect 126020 464176 126026 464188
rect 192662 464176 192668 464188
rect 192720 464176 192726 464228
rect 138474 464108 138480 464160
rect 138532 464148 138538 464160
rect 188614 464148 188620 464160
rect 138532 464120 188620 464148
rect 138532 464108 138538 464120
rect 188614 464108 188620 464120
rect 188672 464108 188678 464160
rect 186682 462952 186688 463004
rect 186740 462992 186746 463004
rect 237466 462992 237472 463004
rect 186740 462964 237472 462992
rect 186740 462952 186746 462964
rect 237466 462952 237472 462964
rect 237524 462952 237530 463004
rect 215938 462340 215944 462392
rect 215996 462380 216002 462392
rect 237374 462380 237380 462392
rect 215996 462352 237380 462380
rect 215996 462340 216002 462352
rect 237374 462340 237380 462352
rect 237432 462340 237438 462392
rect 189074 458260 189080 458312
rect 189132 458300 189138 458312
rect 195238 458300 195244 458312
rect 189132 458272 195244 458300
rect 189132 458260 189138 458272
rect 195238 458260 195244 458272
rect 195296 458260 195302 458312
rect 188430 458192 188436 458244
rect 188488 458232 188494 458244
rect 237374 458232 237380 458244
rect 188488 458204 237380 458232
rect 188488 458192 188494 458204
rect 237374 458192 237380 458204
rect 237432 458192 237438 458244
rect 187234 449828 187240 449880
rect 187292 449868 187298 449880
rect 237374 449868 237380 449880
rect 187292 449840 237380 449868
rect 187292 449828 187298 449840
rect 237374 449828 237380 449840
rect 237432 449828 237438 449880
rect 3326 448536 3332 448588
rect 3384 448576 3390 448588
rect 46198 448576 46204 448588
rect 3384 448548 46204 448576
rect 3384 448536 3390 448548
rect 46198 448536 46204 448548
rect 46256 448536 46262 448588
rect 188522 447108 188528 447160
rect 188580 447148 188586 447160
rect 237374 447148 237380 447160
rect 188580 447120 237380 447148
rect 188580 447108 188586 447120
rect 237374 447108 237380 447120
rect 237432 447108 237438 447160
rect 188614 444320 188620 444372
rect 188672 444360 188678 444372
rect 237374 444360 237380 444372
rect 188672 444332 237380 444360
rect 188672 444320 188678 444332
rect 237374 444320 237380 444332
rect 237432 444320 237438 444372
rect 188614 441600 188620 441652
rect 188672 441640 188678 441652
rect 237374 441640 237380 441652
rect 188672 441612 237380 441640
rect 188672 441600 188678 441612
rect 237374 441600 237380 441612
rect 237432 441600 237438 441652
rect 187142 440172 187148 440224
rect 187200 440212 187206 440224
rect 237374 440212 237380 440224
rect 187200 440184 237380 440212
rect 187200 440172 187206 440184
rect 237374 440172 237380 440184
rect 237432 440172 237438 440224
rect 188706 437452 188712 437504
rect 188764 437492 188770 437504
rect 237374 437492 237380 437504
rect 188764 437464 237380 437492
rect 188764 437452 188770 437464
rect 237374 437452 237380 437464
rect 237432 437452 237438 437504
rect 188798 431944 188804 431996
rect 188856 431984 188862 431996
rect 237374 431984 237380 431996
rect 188856 431956 237380 431984
rect 188856 431944 188862 431956
rect 237374 431944 237380 431956
rect 237432 431944 237438 431996
rect 189994 430584 190000 430636
rect 190052 430624 190058 430636
rect 237374 430624 237380 430636
rect 190052 430596 237380 430624
rect 190052 430584 190058 430596
rect 237374 430584 237380 430596
rect 237432 430584 237438 430636
rect 193950 426504 193956 426556
rect 194008 426544 194014 426556
rect 237374 426544 237380 426556
rect 194008 426516 237380 426544
rect 194008 426504 194014 426516
rect 237374 426504 237380 426516
rect 237432 426504 237438 426556
rect 188890 426436 188896 426488
rect 188948 426476 188954 426488
rect 237466 426476 237472 426488
rect 188948 426448 237472 426476
rect 188948 426436 188954 426448
rect 237466 426436 237472 426448
rect 237524 426436 237530 426488
rect 187050 423580 187056 423632
rect 187108 423620 187114 423632
rect 237374 423620 237380 423632
rect 187108 423592 237380 423620
rect 187108 423580 187114 423592
rect 237374 423580 237380 423592
rect 237432 423580 237438 423632
rect 188982 422288 188988 422340
rect 189040 422328 189046 422340
rect 237374 422328 237380 422340
rect 189040 422300 237380 422328
rect 189040 422288 189046 422300
rect 237374 422288 237380 422300
rect 237432 422288 237438 422340
rect 192662 419432 192668 419484
rect 192720 419472 192726 419484
rect 237374 419472 237380 419484
rect 192720 419444 237380 419472
rect 192720 419432 192726 419444
rect 237374 419432 237380 419444
rect 237432 419432 237438 419484
rect 538950 418140 538956 418192
rect 539008 418180 539014 418192
rect 579614 418180 579620 418192
rect 539008 418152 579620 418180
rect 539008 418140 539014 418152
rect 579614 418140 579620 418152
rect 579672 418140 579678 418192
rect 187050 416780 187056 416832
rect 187108 416820 187114 416832
rect 237374 416820 237380 416832
rect 187108 416792 237380 416820
rect 187108 416780 187114 416792
rect 237374 416780 237380 416792
rect 237432 416780 237438 416832
rect 187142 415420 187148 415472
rect 187200 415460 187206 415472
rect 237374 415460 237380 415472
rect 187200 415432 237380 415460
rect 187200 415420 187206 415432
rect 237374 415420 237380 415432
rect 237432 415420 237438 415472
rect 190086 413924 190092 413976
rect 190144 413964 190150 413976
rect 237374 413964 237380 413976
rect 190144 413936 237380 413964
rect 190144 413924 190150 413936
rect 237374 413924 237380 413936
rect 237432 413924 237438 413976
rect 187234 411272 187240 411324
rect 187292 411312 187298 411324
rect 237374 411312 237380 411324
rect 187292 411284 237380 411312
rect 187292 411272 187298 411284
rect 237374 411272 237380 411284
rect 237432 411272 237438 411324
rect 189902 408416 189908 408468
rect 189960 408456 189966 408468
rect 237374 408456 237380 408468
rect 189960 408428 237380 408456
rect 189960 408416 189966 408428
rect 237374 408416 237380 408428
rect 237432 408416 237438 408468
rect 189902 405696 189908 405748
rect 189960 405736 189966 405748
rect 237374 405736 237380 405748
rect 189960 405708 237380 405736
rect 189960 405696 189966 405708
rect 237374 405696 237380 405708
rect 237432 405696 237438 405748
rect 187326 401616 187332 401668
rect 187384 401656 187390 401668
rect 237374 401656 237380 401668
rect 187384 401628 237380 401656
rect 187384 401616 187390 401628
rect 237374 401616 237380 401628
rect 237432 401616 237438 401668
rect 190086 400188 190092 400240
rect 190144 400228 190150 400240
rect 237374 400228 237380 400240
rect 190144 400200 237380 400228
rect 190144 400188 190150 400200
rect 237374 400188 237380 400200
rect 237432 400188 237438 400240
rect 189074 398828 189080 398880
rect 189132 398868 189138 398880
rect 192662 398868 192668 398880
rect 189132 398840 192668 398868
rect 189132 398828 189138 398840
rect 192662 398828 192668 398840
rect 192720 398828 192726 398880
rect 3326 397468 3332 397520
rect 3384 397508 3390 397520
rect 44818 397508 44824 397520
rect 3384 397480 44824 397508
rect 3384 397468 3390 397480
rect 44818 397468 44824 397480
rect 44876 397468 44882 397520
rect 189074 397468 189080 397520
rect 189132 397508 189138 397520
rect 192754 397508 192760 397520
rect 189132 397480 192760 397508
rect 189132 397468 189138 397480
rect 192754 397468 192760 397480
rect 192812 397468 192818 397520
rect 189074 396176 189080 396228
rect 189132 396216 189138 396228
rect 195330 396216 195336 396228
rect 189132 396188 195336 396216
rect 189132 396176 189138 396188
rect 195330 396176 195336 396188
rect 195388 396176 195394 396228
rect 190178 396108 190184 396160
rect 190236 396148 190242 396160
rect 237374 396148 237380 396160
rect 190236 396120 237380 396148
rect 190236 396108 190242 396120
rect 237374 396108 237380 396120
rect 237432 396108 237438 396160
rect 187418 396040 187424 396092
rect 187476 396080 187482 396092
rect 237466 396080 237472 396092
rect 187476 396052 237472 396080
rect 187476 396040 187482 396052
rect 237466 396040 237472 396052
rect 237524 396040 237530 396092
rect 189442 394680 189448 394732
rect 189500 394720 189506 394732
rect 195422 394720 195428 394732
rect 189500 394692 195428 394720
rect 189500 394680 189506 394692
rect 195422 394680 195428 394692
rect 195480 394680 195486 394732
rect 189074 393320 189080 393372
rect 189132 393360 189138 393372
rect 195514 393360 195520 393372
rect 189132 393332 195520 393360
rect 189132 393320 189138 393332
rect 195514 393320 195520 393332
rect 195572 393320 195578 393372
rect 187510 391960 187516 392012
rect 187568 392000 187574 392012
rect 237374 392000 237380 392012
rect 187568 391972 237380 392000
rect 187568 391960 187574 391972
rect 237374 391960 237380 391972
rect 237432 391960 237438 392012
rect 188246 390532 188252 390584
rect 188304 390572 188310 390584
rect 237374 390572 237380 390584
rect 188304 390544 237380 390572
rect 188304 390532 188310 390544
rect 237374 390532 237380 390544
rect 237432 390532 237438 390584
rect 186958 389104 186964 389156
rect 187016 389144 187022 389156
rect 237374 389144 237380 389156
rect 187016 389116 237380 389144
rect 187016 389104 187022 389116
rect 237374 389104 237380 389116
rect 237432 389104 237438 389156
rect 186958 386384 186964 386436
rect 187016 386424 187022 386436
rect 237374 386424 237380 386436
rect 187016 386396 237380 386424
rect 187016 386384 187022 386396
rect 237374 386384 237380 386396
rect 237432 386384 237438 386436
rect 187786 385024 187792 385076
rect 187844 385064 187850 385076
rect 237374 385064 237380 385076
rect 187844 385036 237380 385064
rect 187844 385024 187850 385036
rect 237374 385024 237380 385036
rect 237432 385024 237438 385076
rect 188338 383596 188344 383648
rect 188396 383636 188402 383648
rect 237374 383636 237380 383648
rect 188396 383608 237380 383636
rect 188396 383596 188402 383608
rect 237374 383596 237380 383608
rect 237432 383596 237438 383648
rect 187694 380876 187700 380928
rect 187752 380916 187758 380928
rect 237374 380916 237380 380928
rect 187752 380888 237380 380916
rect 187752 380876 187758 380888
rect 237374 380876 237380 380888
rect 237432 380876 237438 380928
rect 186682 380128 186688 380180
rect 186740 380168 186746 380180
rect 237926 380168 237932 380180
rect 186740 380140 237932 380168
rect 186740 380128 186746 380140
rect 237926 380128 237932 380140
rect 237984 380128 237990 380180
rect 48222 379516 48228 379568
rect 48280 379556 48286 379568
rect 49878 379556 49884 379568
rect 48280 379528 49884 379556
rect 48280 379516 48286 379528
rect 49878 379516 49884 379528
rect 49936 379516 49942 379568
rect 116026 379448 116032 379500
rect 116084 379488 116090 379500
rect 187418 379488 187424 379500
rect 116084 379460 187424 379488
rect 116084 379448 116090 379460
rect 187418 379448 187424 379460
rect 187476 379448 187482 379500
rect 113542 379380 113548 379432
rect 113600 379420 113606 379432
rect 187510 379420 187516 379432
rect 113600 379392 187516 379420
rect 113600 379380 113606 379392
rect 187510 379380 187516 379392
rect 187568 379380 187574 379432
rect 110966 379312 110972 379364
rect 111024 379352 111030 379364
rect 186958 379352 186964 379364
rect 111024 379324 186964 379352
rect 111024 379312 111030 379324
rect 186958 379312 186964 379324
rect 187016 379312 187022 379364
rect 150986 379244 150992 379296
rect 151044 379284 151050 379296
rect 235902 379284 235908 379296
rect 151044 379256 235908 379284
rect 151044 379244 151050 379256
rect 235902 379244 235908 379256
rect 235960 379244 235966 379296
rect 144914 379176 144920 379228
rect 144972 379216 144978 379228
rect 238018 379216 238024 379228
rect 144972 379188 238024 379216
rect 144972 379176 144978 379188
rect 238018 379176 238024 379188
rect 238076 379176 238082 379228
rect 89438 379108 89444 379160
rect 89496 379148 89502 379160
rect 188246 379148 188252 379160
rect 89496 379120 188252 379148
rect 89496 379108 89502 379120
rect 188246 379108 188252 379120
rect 188304 379108 188310 379160
rect 88150 379040 88156 379092
rect 88208 379080 88214 379092
rect 187786 379080 187792 379092
rect 88208 379052 187792 379080
rect 88208 379040 88214 379052
rect 187786 379040 187792 379052
rect 187844 379040 187850 379092
rect 90726 378972 90732 379024
rect 90784 379012 90790 379024
rect 190178 379012 190184 379024
rect 90784 378984 190184 379012
rect 90784 378972 90790 378984
rect 190178 378972 190184 378984
rect 190236 378972 190242 379024
rect 87046 378904 87052 378956
rect 87104 378944 87110 378956
rect 187694 378944 187700 378956
rect 87104 378916 187700 378944
rect 87104 378904 87110 378916
rect 187694 378904 187700 378916
rect 187752 378904 187758 378956
rect 135990 378836 135996 378888
rect 136048 378876 136054 378888
rect 237466 378876 237472 378888
rect 136048 378848 237472 378876
rect 136048 378836 136054 378848
rect 237466 378836 237472 378848
rect 237524 378836 237530 378888
rect 120994 378768 121000 378820
rect 121052 378808 121058 378820
rect 237834 378808 237840 378820
rect 121052 378780 237840 378808
rect 121052 378768 121058 378780
rect 237834 378768 237840 378780
rect 237892 378768 237898 378820
rect 118326 378700 118332 378752
rect 118384 378740 118390 378752
rect 187326 378740 187332 378752
rect 118384 378712 187332 378740
rect 118384 378700 118390 378712
rect 187326 378700 187332 378712
rect 187384 378700 187390 378752
rect 123478 378632 123484 378684
rect 123536 378672 123542 378684
rect 187234 378672 187240 378684
rect 123536 378644 187240 378672
rect 123536 378632 123542 378644
rect 187234 378632 187240 378644
rect 187292 378632 187298 378684
rect 130930 378564 130936 378616
rect 130988 378604 130994 378616
rect 188890 378604 188896 378616
rect 130988 378576 188896 378604
rect 130988 378564 130994 378576
rect 188890 378564 188896 378576
rect 188948 378564 188954 378616
rect 542998 378156 543004 378208
rect 543056 378196 543062 378208
rect 580166 378196 580172 378208
rect 543056 378168 580172 378196
rect 543056 378156 543062 378168
rect 580166 378156 580172 378168
rect 580224 378156 580230 378208
rect 91922 378020 91928 378072
rect 91980 378060 91986 378072
rect 190086 378060 190092 378072
rect 91980 378032 190092 378060
rect 91980 378020 91986 378032
rect 190086 378020 190092 378032
rect 190144 378020 190150 378072
rect 198182 378020 198188 378072
rect 198240 378060 198246 378072
rect 237374 378060 237380 378072
rect 198240 378032 237380 378060
rect 198240 378020 198246 378032
rect 237374 378020 237380 378032
rect 237432 378020 237438 378072
rect 92842 377952 92848 378004
rect 92900 377992 92906 378004
rect 189902 377992 189908 378004
rect 92900 377964 189908 377992
rect 92900 377952 92906 377964
rect 189902 377952 189908 377964
rect 189960 377952 189966 378004
rect 93946 377884 93952 377936
rect 94004 377924 94010 377936
rect 186682 377924 186688 377936
rect 94004 377896 186688 377924
rect 94004 377884 94010 377896
rect 186682 377884 186688 377896
rect 186740 377884 186746 377936
rect 95234 377816 95240 377868
rect 95292 377856 95298 377868
rect 187142 377856 187148 377868
rect 95292 377828 187148 377856
rect 95292 377816 95298 377828
rect 187142 377816 187148 377828
rect 187200 377816 187206 377868
rect 96430 377748 96436 377800
rect 96488 377788 96494 377800
rect 140774 377788 140780 377800
rect 96488 377760 140780 377788
rect 96488 377748 96494 377760
rect 140774 377748 140780 377760
rect 140832 377748 140838 377800
rect 148594 377748 148600 377800
rect 148652 377788 148658 377800
rect 215938 377788 215944 377800
rect 148652 377760 215944 377788
rect 148652 377748 148658 377760
rect 215938 377748 215944 377760
rect 215996 377748 216002 377800
rect 125962 377680 125968 377732
rect 126020 377720 126026 377732
rect 187050 377720 187056 377732
rect 126020 377692 187056 377720
rect 126020 377680 126026 377692
rect 187050 377680 187056 377692
rect 187108 377680 187114 377732
rect 128538 377612 128544 377664
rect 128596 377652 128602 377664
rect 188982 377652 188988 377664
rect 128596 377624 188988 377652
rect 128596 377612 128602 377624
rect 188982 377612 188988 377624
rect 189040 377612 189046 377664
rect 133506 377544 133512 377596
rect 133564 377584 133570 377596
rect 188798 377584 188804 377596
rect 133564 377556 188804 377584
rect 133564 377544 133570 377556
rect 188798 377544 188804 377556
rect 188856 377544 188862 377596
rect 108482 377476 108488 377528
rect 108540 377516 108546 377528
rect 135990 377516 135996 377528
rect 108540 377488 135996 377516
rect 108540 377476 108546 377488
rect 135990 377476 135996 377488
rect 136048 377476 136054 377528
rect 136082 377476 136088 377528
rect 136140 377516 136146 377528
rect 188706 377516 188712 377528
rect 136140 377488 188712 377516
rect 136140 377476 136146 377488
rect 188706 377476 188712 377488
rect 188764 377476 188770 377528
rect 106090 377408 106096 377460
rect 106148 377448 106154 377460
rect 237374 377448 237380 377460
rect 106148 377420 237380 377448
rect 106148 377408 106154 377420
rect 237374 377408 237380 377420
rect 237432 377408 237438 377460
rect 138658 377340 138664 377392
rect 138716 377380 138722 377392
rect 188614 377380 188620 377392
rect 138716 377352 188620 377380
rect 138716 377340 138722 377352
rect 188614 377340 188620 377352
rect 188672 377340 188678 377392
rect 141142 377272 141148 377324
rect 141200 377312 141206 377324
rect 188522 377312 188528 377324
rect 141200 377284 188528 377312
rect 141200 377272 141206 377284
rect 188522 377272 188528 377284
rect 188580 377272 188586 377324
rect 146018 377204 146024 377256
rect 146076 377244 146082 377256
rect 188430 377244 188436 377256
rect 146076 377216 188436 377244
rect 146076 377204 146082 377216
rect 188430 377204 188436 377216
rect 188488 377204 188494 377256
rect 99926 377136 99932 377188
rect 99984 377176 99990 377188
rect 238570 377176 238576 377188
rect 99984 377148 238576 377176
rect 99984 377136 99990 377148
rect 238570 377136 238576 377148
rect 238628 377136 238634 377188
rect 78306 377000 78312 377052
rect 78364 377040 78370 377052
rect 79318 377040 79324 377052
rect 78364 377012 79324 377040
rect 78364 377000 78370 377012
rect 79318 377000 79324 377012
rect 79376 377000 79382 377052
rect 85942 376660 85948 376712
rect 86000 376700 86006 376712
rect 237374 376700 237380 376712
rect 86000 376672 237380 376700
rect 86000 376660 86006 376672
rect 237374 376660 237380 376672
rect 237432 376660 237438 376712
rect 97626 376592 97632 376644
rect 97684 376632 97690 376644
rect 193950 376632 193956 376644
rect 97684 376604 193956 376632
rect 97684 376592 97690 376604
rect 193950 376592 193956 376604
rect 194008 376592 194014 376644
rect 153378 376524 153384 376576
rect 153436 376564 153442 376576
rect 235718 376564 235724 376576
rect 153436 376536 235724 376564
rect 153436 376524 153442 376536
rect 235718 376524 235724 376536
rect 235776 376524 235782 376576
rect 155954 376456 155960 376508
rect 156012 376496 156018 376508
rect 235534 376496 235540 376508
rect 156012 376468 235540 376496
rect 156012 376456 156018 376468
rect 235534 376456 235540 376468
rect 235592 376456 235598 376508
rect 49326 375980 49332 376032
rect 49384 376020 49390 376032
rect 238018 376020 238024 376032
rect 49384 375992 238024 376020
rect 49384 375980 49390 375992
rect 238018 375980 238024 375992
rect 238076 375980 238082 376032
rect 198090 373940 198096 373992
rect 198148 373980 198154 373992
rect 237374 373980 237380 373992
rect 198148 373952 237380 373980
rect 198148 373940 198154 373952
rect 237374 373940 237380 373952
rect 237432 373940 237438 373992
rect 104802 372512 104808 372564
rect 104860 372552 104866 372564
rect 237374 372552 237380 372564
rect 104860 372524 237380 372552
rect 104860 372512 104866 372524
rect 237374 372512 237380 372524
rect 237432 372512 237438 372564
rect 47854 371832 47860 371884
rect 47912 371872 47918 371884
rect 122098 371872 122104 371884
rect 47912 371844 122104 371872
rect 47912 371832 47918 371844
rect 122098 371832 122104 371844
rect 122156 371832 122162 371884
rect 85482 371152 85488 371204
rect 85540 371192 85546 371204
rect 237374 371192 237380 371204
rect 85540 371164 237380 371192
rect 85540 371152 85546 371164
rect 237374 371152 237380 371164
rect 237432 371152 237438 371204
rect 47946 369112 47952 369164
rect 48004 369152 48010 369164
rect 177298 369152 177304 369164
rect 48004 369124 177304 369152
rect 48004 369112 48010 369124
rect 177298 369112 177304 369124
rect 177356 369112 177362 369164
rect 191282 368432 191288 368484
rect 191340 368472 191346 368484
rect 237374 368472 237380 368484
rect 191340 368444 237380 368472
rect 191340 368432 191346 368444
rect 237374 368432 237380 368444
rect 237432 368432 237438 368484
rect 84010 367004 84016 367056
rect 84068 367044 84074 367056
rect 237466 367044 237472 367056
rect 84068 367016 237472 367044
rect 84068 367004 84074 367016
rect 237466 367004 237472 367016
rect 237524 367004 237530 367056
rect 102042 366936 102048 366988
rect 102100 366976 102106 366988
rect 237374 366976 237380 366988
rect 102100 366948 237380 366976
rect 102100 366936 102106 366948
rect 237374 366936 237380 366948
rect 237432 366936 237438 366988
rect 49418 364964 49424 365016
rect 49476 365004 49482 365016
rect 238110 365004 238116 365016
rect 49476 364976 238116 365004
rect 49476 364964 49482 364976
rect 238110 364964 238116 364976
rect 238168 364964 238174 365016
rect 538950 364352 538956 364404
rect 539008 364392 539014 364404
rect 580166 364392 580172 364404
rect 539008 364364 580172 364392
rect 539008 364352 539014 364364
rect 580166 364352 580172 364364
rect 580224 364352 580230 364404
rect 99282 362856 99288 362908
rect 99340 362896 99346 362908
rect 237466 362896 237472 362908
rect 99340 362868 237472 362896
rect 99340 362856 99346 362868
rect 237466 362856 237472 362868
rect 237524 362856 237530 362908
rect 199378 362788 199384 362840
rect 199436 362828 199442 362840
rect 237374 362828 237380 362840
rect 199436 362800 237380 362828
rect 199436 362788 199442 362800
rect 237374 362788 237380 362800
rect 237432 362788 237438 362840
rect 82722 361496 82728 361548
rect 82780 361536 82786 361548
rect 237374 361536 237380 361548
rect 82780 361508 237380 361536
rect 82780 361496 82786 361508
rect 237374 361496 237380 361508
rect 237432 361496 237438 361548
rect 173710 360136 173716 360188
rect 173768 360176 173774 360188
rect 237374 360176 237380 360188
rect 173768 360148 237380 360176
rect 173768 360136 173774 360148
rect 237374 360136 237380 360148
rect 237432 360136 237438 360188
rect 48038 358708 48044 358760
rect 48096 358748 48102 358760
rect 237374 358748 237380 358760
rect 48096 358720 237380 358748
rect 48096 358708 48102 358720
rect 237374 358708 237380 358720
rect 237432 358708 237438 358760
rect 191190 358640 191196 358692
rect 191248 358680 191254 358692
rect 237466 358680 237472 358692
rect 191248 358652 237472 358680
rect 191248 358640 191254 358652
rect 237466 358640 237472 358652
rect 237524 358640 237530 358692
rect 96522 357348 96528 357400
rect 96580 357388 96586 357400
rect 237374 357388 237380 357400
rect 96580 357360 237380 357388
rect 96580 357348 96586 357360
rect 237374 357348 237380 357360
rect 237432 357348 237438 357400
rect 81158 355988 81164 356040
rect 81216 356028 81222 356040
rect 237374 356028 237380 356040
rect 81216 356000 237380 356028
rect 81216 355988 81222 356000
rect 237374 355988 237380 356000
rect 237432 355988 237438 356040
rect 173802 355920 173808 355972
rect 173860 355960 173866 355972
rect 237466 355960 237472 355972
rect 173860 355932 237472 355960
rect 173860 355920 173866 355932
rect 237466 355920 237472 355932
rect 237524 355920 237530 355972
rect 177298 354628 177304 354680
rect 177356 354668 177362 354680
rect 237374 354668 237380 354680
rect 177356 354640 237380 354668
rect 177356 354628 177362 354640
rect 237374 354628 237380 354640
rect 237432 354628 237438 354680
rect 197998 353200 198004 353252
rect 198056 353240 198062 353252
rect 237374 353240 237380 353252
rect 198056 353212 237380 353240
rect 198056 353200 198062 353212
rect 237374 353200 237380 353212
rect 237432 353200 237438 353252
rect 81250 351840 81256 351892
rect 81308 351880 81314 351892
rect 237466 351880 237472 351892
rect 81308 351852 237472 351880
rect 81308 351840 81314 351852
rect 237466 351840 237472 351852
rect 237524 351840 237530 351892
rect 93762 351772 93768 351824
rect 93820 351812 93826 351824
rect 237374 351812 237380 351824
rect 93820 351784 237380 351812
rect 93820 351772 93826 351784
rect 237374 351772 237380 351784
rect 237432 351772 237438 351824
rect 195514 350480 195520 350532
rect 195572 350520 195578 350532
rect 237374 350520 237380 350532
rect 195572 350492 237380 350520
rect 195572 350480 195578 350492
rect 237374 350480 237380 350492
rect 237432 350480 237438 350532
rect 49878 349052 49884 349104
rect 49936 349092 49942 349104
rect 237374 349092 237380 349104
rect 49936 349064 237380 349092
rect 49936 349052 49942 349064
rect 237374 349052 237380 349064
rect 237432 349052 237438 349104
rect 92382 347692 92388 347744
rect 92440 347732 92446 347744
rect 237374 347732 237380 347744
rect 92440 347704 237380 347732
rect 92440 347692 92446 347704
rect 237374 347692 237380 347704
rect 237432 347692 237438 347744
rect 235442 347624 235448 347676
rect 235500 347664 235506 347676
rect 237466 347664 237472 347676
rect 235500 347636 237472 347664
rect 235500 347624 235506 347636
rect 237466 347624 237472 347636
rect 237524 347624 237530 347676
rect 79962 346332 79968 346384
rect 80020 346372 80026 346384
rect 237374 346372 237380 346384
rect 80020 346344 237380 346372
rect 80020 346332 80026 346344
rect 237374 346332 237380 346344
rect 237432 346332 237438 346384
rect 3050 345040 3056 345092
rect 3108 345080 3114 345092
rect 233878 345080 233884 345092
rect 3108 345052 233884 345080
rect 3108 345040 3114 345052
rect 233878 345040 233884 345052
rect 233936 345040 233942 345092
rect 195422 344972 195428 345024
rect 195480 345012 195486 345024
rect 237374 345012 237380 345024
rect 195480 344984 237380 345012
rect 195480 344972 195486 344984
rect 237374 344972 237380 344984
rect 237432 344972 237438 345024
rect 196618 343544 196624 343596
rect 196676 343584 196682 343596
rect 237374 343584 237380 343596
rect 196676 343556 237380 343584
rect 196676 343544 196682 343556
rect 237374 343544 237380 343556
rect 237432 343544 237438 343596
rect 89622 342184 89628 342236
rect 89680 342224 89686 342236
rect 237374 342224 237380 342236
rect 89680 342196 237380 342224
rect 89680 342184 89686 342196
rect 237374 342184 237380 342196
rect 237432 342184 237438 342236
rect 78490 340824 78496 340876
rect 78548 340864 78554 340876
rect 237374 340864 237380 340876
rect 78548 340836 237380 340864
rect 78548 340824 78554 340836
rect 237374 340824 237380 340836
rect 237432 340824 237438 340876
rect 195330 340756 195336 340808
rect 195388 340796 195394 340808
rect 237466 340796 237472 340808
rect 195388 340768 237472 340796
rect 195388 340756 195394 340768
rect 237466 340756 237472 340768
rect 237524 340756 237530 340808
rect 73062 338036 73068 338088
rect 73120 338076 73126 338088
rect 237374 338076 237380 338088
rect 73120 338048 237380 338076
rect 73120 338036 73126 338048
rect 237374 338036 237380 338048
rect 237432 338036 237438 338088
rect 86770 336676 86776 336728
rect 86828 336716 86834 336728
rect 237466 336716 237472 336728
rect 86828 336688 237472 336716
rect 86828 336676 86834 336688
rect 237466 336676 237472 336688
rect 237524 336676 237530 336728
rect 189810 336608 189816 336660
rect 189868 336648 189874 336660
rect 237374 336648 237380 336660
rect 189868 336620 237380 336648
rect 189868 336608 189874 336620
rect 237374 336608 237380 336620
rect 237432 336608 237438 336660
rect 77202 335248 77208 335300
rect 77260 335288 77266 335300
rect 237374 335288 237380 335300
rect 77260 335260 237380 335288
rect 77260 335248 77266 335260
rect 237374 335248 237380 335260
rect 237432 335248 237438 335300
rect 192754 333888 192760 333940
rect 192812 333928 192818 333940
rect 237374 333928 237380 333940
rect 192812 333900 237380 333928
rect 192812 333888 192818 333900
rect 237374 333888 237380 333900
rect 237432 333888 237438 333940
rect 49234 332528 49240 332580
rect 49292 332568 49298 332580
rect 237374 332568 237380 332580
rect 49292 332540 237380 332568
rect 49292 332528 49298 332540
rect 237374 332528 237380 332540
rect 237432 332528 237438 332580
rect 71682 332460 71688 332512
rect 71740 332500 71746 332512
rect 237466 332500 237472 332512
rect 71740 332472 237472 332500
rect 71740 332460 71746 332472
rect 237466 332460 237472 332472
rect 237524 332460 237530 332512
rect 193858 331168 193864 331220
rect 193916 331208 193922 331220
rect 237374 331208 237380 331220
rect 193916 331180 237380 331208
rect 193916 331168 193922 331180
rect 237374 331168 237380 331180
rect 237432 331168 237438 331220
rect 75822 329740 75828 329792
rect 75880 329780 75886 329792
rect 237466 329780 237472 329792
rect 75880 329752 237472 329780
rect 75880 329740 75886 329752
rect 237466 329740 237472 329752
rect 237524 329740 237530 329792
rect 84102 329672 84108 329724
rect 84160 329712 84166 329724
rect 237374 329712 237380 329724
rect 84160 329684 237380 329712
rect 84160 329672 84166 329684
rect 237374 329672 237380 329684
rect 237432 329672 237438 329724
rect 192662 328380 192668 328432
rect 192720 328420 192726 328432
rect 237374 328420 237380 328432
rect 192720 328392 237380 328420
rect 192720 328380 192726 328392
rect 237374 328380 237380 328392
rect 237432 328380 237438 328432
rect 49602 327020 49608 327072
rect 49660 327060 49666 327072
rect 237374 327060 237380 327072
rect 49660 327032 237380 327060
rect 49660 327020 49666 327032
rect 237374 327020 237380 327032
rect 237432 327020 237438 327072
rect 70302 325592 70308 325644
rect 70360 325632 70366 325644
rect 237374 325632 237380 325644
rect 70360 325604 237380 325632
rect 70360 325592 70366 325604
rect 237374 325592 237380 325604
rect 237432 325592 237438 325644
rect 235350 325320 235356 325372
rect 235408 325360 235414 325372
rect 237374 325360 237380 325372
rect 235408 325332 237380 325360
rect 235408 325320 235414 325332
rect 237374 325320 237380 325332
rect 237432 325320 237438 325372
rect 74350 324912 74356 324964
rect 74408 324952 74414 324964
rect 237466 324952 237472 324964
rect 74408 324924 237472 324952
rect 74408 324912 74414 324924
rect 237466 324912 237472 324924
rect 237524 324912 237530 324964
rect 540238 324300 540244 324352
rect 540296 324340 540302 324352
rect 579614 324340 579620 324352
rect 540296 324312 579620 324340
rect 540296 324300 540302 324312
rect 579614 324300 579620 324312
rect 579672 324300 579678 324352
rect 81342 324232 81348 324284
rect 81400 324272 81406 324284
rect 237374 324272 237380 324284
rect 81400 324244 237380 324272
rect 81400 324232 81406 324244
rect 237374 324232 237380 324244
rect 237432 324232 237438 324284
rect 74442 323552 74448 323604
rect 74500 323592 74506 323604
rect 237558 323592 237564 323604
rect 74500 323564 237564 323592
rect 74500 323552 74506 323564
rect 237558 323552 237564 323564
rect 237616 323552 237622 323604
rect 67542 321512 67548 321564
rect 67600 321552 67606 321564
rect 237466 321552 237472 321564
rect 67600 321524 237472 321552
rect 67600 321512 67606 321524
rect 237466 321512 237472 321524
rect 237524 321512 237530 321564
rect 192570 321444 192576 321496
rect 192628 321484 192634 321496
rect 237374 321484 237380 321496
rect 192628 321456 237380 321484
rect 192628 321444 192634 321456
rect 237374 321444 237380 321456
rect 237432 321444 237438 321496
rect 68922 320084 68928 320136
rect 68980 320124 68986 320136
rect 237374 320124 237380 320136
rect 68980 320096 237380 320124
rect 68980 320084 68986 320096
rect 237374 320084 237380 320096
rect 237432 320084 237438 320136
rect 79318 317364 79324 317416
rect 79376 317404 79382 317416
rect 237374 317404 237380 317416
rect 79376 317376 237380 317404
rect 79376 317364 79382 317376
rect 237374 317364 237380 317376
rect 237432 317364 237438 317416
rect 192478 315936 192484 315988
rect 192536 315976 192542 315988
rect 237374 315976 237380 315988
rect 192536 315948 237380 315976
rect 192536 315936 192542 315948
rect 237374 315936 237380 315948
rect 237432 315936 237438 315988
rect 66162 314576 66168 314628
rect 66220 314616 66226 314628
rect 237374 314616 237380 314628
rect 66220 314588 237380 314616
rect 66220 314576 66226 314588
rect 237374 314576 237380 314588
rect 237432 314576 237438 314628
rect 48130 313216 48136 313268
rect 48188 313256 48194 313268
rect 237374 313256 237380 313268
rect 48188 313228 237380 313256
rect 48188 313216 48194 313228
rect 237374 313216 237380 313228
rect 237432 313216 237438 313268
rect 195238 313148 195244 313200
rect 195296 313188 195302 313200
rect 237466 313188 237472 313200
rect 195296 313160 237472 313188
rect 195296 313148 195302 313160
rect 237466 313148 237472 313160
rect 237524 313148 237530 313200
rect 122098 311788 122104 311840
rect 122156 311828 122162 311840
rect 237374 311828 237380 311840
rect 122156 311800 237380 311828
rect 122156 311788 122162 311800
rect 237374 311788 237380 311800
rect 237432 311788 237438 311840
rect 232498 309204 232504 309256
rect 232556 309244 232562 309256
rect 237466 309244 237472 309256
rect 232556 309216 237472 309244
rect 232556 309204 232562 309216
rect 237466 309204 237472 309216
rect 237524 309204 237530 309256
rect 157242 309136 157248 309188
rect 157300 309176 157306 309188
rect 237374 309176 237380 309188
rect 157300 309148 237380 309176
rect 157300 309136 157306 309148
rect 237374 309136 237380 309148
rect 237432 309136 237438 309188
rect 235350 307776 235356 307828
rect 235408 307816 235414 307828
rect 237374 307816 237380 307828
rect 235408 307788 237380 307816
rect 235408 307776 235414 307788
rect 237374 307776 237380 307788
rect 237432 307776 237438 307828
rect 232590 305056 232596 305108
rect 232648 305096 232654 305108
rect 237466 305096 237472 305108
rect 232648 305068 237472 305096
rect 232648 305056 232654 305068
rect 237466 305056 237472 305068
rect 237524 305056 237530 305108
rect 235442 304988 235448 305040
rect 235500 305028 235506 305040
rect 237374 305028 237380 305040
rect 235500 305000 237380 305028
rect 235500 304988 235506 305000
rect 237374 304988 237380 305000
rect 237432 304988 237438 305040
rect 151722 303628 151728 303680
rect 151780 303668 151786 303680
rect 237374 303668 237380 303680
rect 151780 303640 237380 303668
rect 151780 303628 151786 303640
rect 237374 303628 237380 303640
rect 237432 303628 237438 303680
rect 232682 302200 232688 302252
rect 232740 302240 232746 302252
rect 237374 302240 237380 302252
rect 232740 302212 237380 302240
rect 232740 302200 232746 302212
rect 237374 302200 237380 302212
rect 237432 302200 237438 302252
rect 235534 300908 235540 300960
rect 235592 300948 235598 300960
rect 237466 300948 237472 300960
rect 235592 300920 237472 300948
rect 235592 300908 235598 300920
rect 237466 300908 237472 300920
rect 237524 300908 237530 300960
rect 148962 300840 148968 300892
rect 149020 300880 149026 300892
rect 237374 300880 237380 300892
rect 149020 300852 237380 300880
rect 149020 300840 149026 300852
rect 237374 300840 237380 300852
rect 237432 300840 237438 300892
rect 235626 298120 235632 298172
rect 235684 298160 235690 298172
rect 237374 298160 237380 298172
rect 235684 298132 237380 298160
rect 235684 298120 235690 298132
rect 237374 298120 237380 298132
rect 237432 298120 237438 298172
rect 146202 296692 146208 296744
rect 146260 296732 146266 296744
rect 237374 296732 237380 296744
rect 146260 296704 237380 296732
rect 146260 296692 146266 296704
rect 237374 296692 237380 296704
rect 237432 296692 237438 296744
rect 235718 295332 235724 295384
rect 235776 295372 235782 295384
rect 237374 295372 237380 295384
rect 235776 295344 237380 295372
rect 235776 295332 235782 295344
rect 237374 295332 237380 295344
rect 237432 295332 237438 295384
rect 144822 293972 144828 294024
rect 144880 294012 144886 294024
rect 237374 294012 237380 294024
rect 144880 293984 237380 294012
rect 144880 293972 144886 293984
rect 237374 293972 237380 293984
rect 237432 293972 237438 294024
rect 3142 292612 3148 292664
rect 3200 292652 3206 292664
rect 236638 292652 236644 292664
rect 3200 292624 236644 292652
rect 3200 292612 3206 292624
rect 236638 292612 236644 292624
rect 236696 292612 236702 292664
rect 235902 292544 235908 292596
rect 235960 292584 235966 292596
rect 237374 292584 237380 292596
rect 235960 292556 237380 292584
rect 235960 292544 235966 292556
rect 237374 292544 237380 292556
rect 237432 292544 237438 292596
rect 142062 291184 142068 291236
rect 142120 291224 142126 291236
rect 237374 291224 237380 291236
rect 142120 291196 237380 291224
rect 142120 291184 142126 291196
rect 237374 291184 237380 291196
rect 237432 291184 237438 291236
rect 154482 290436 154488 290488
rect 154540 290476 154546 290488
rect 238018 290476 238024 290488
rect 154540 290448 238024 290476
rect 154540 290436 154546 290448
rect 238018 290436 238024 290448
rect 238076 290436 238082 290488
rect 235166 289824 235172 289876
rect 235224 289864 235230 289876
rect 237374 289864 237380 289876
rect 235224 289836 237380 289864
rect 235224 289824 235230 289836
rect 237374 289824 237380 289836
rect 237432 289824 237438 289876
rect 139302 288396 139308 288448
rect 139360 288436 139366 288448
rect 237374 288436 237380 288448
rect 139360 288408 237380 288436
rect 139360 288396 139366 288408
rect 237374 288396 237380 288408
rect 237432 288396 237438 288448
rect 117222 286492 117228 286544
rect 117280 286532 117286 286544
rect 169754 286532 169760 286544
rect 117280 286504 169760 286532
rect 117280 286492 117286 286504
rect 169754 286492 169760 286504
rect 169812 286492 169818 286544
rect 170674 286492 170680 286544
rect 170732 286532 170738 286544
rect 192478 286532 192484 286544
rect 170732 286504 192484 286532
rect 170732 286492 170738 286504
rect 192478 286492 192484 286504
rect 192536 286492 192542 286544
rect 121362 286424 121368 286476
rect 121420 286464 121426 286476
rect 137278 286464 137284 286476
rect 121420 286436 137284 286464
rect 121420 286424 121426 286436
rect 137278 286424 137284 286436
rect 137336 286424 137342 286476
rect 169662 286424 169668 286476
rect 169720 286464 169726 286476
rect 192662 286464 192668 286476
rect 169720 286436 192668 286464
rect 169720 286424 169726 286436
rect 192662 286424 192668 286436
rect 192720 286424 192726 286476
rect 136542 286356 136548 286408
rect 136600 286396 136606 286408
rect 237374 286396 237380 286408
rect 136600 286368 237380 286396
rect 136600 286356 136606 286368
rect 237374 286356 237380 286368
rect 237432 286356 237438 286408
rect 49602 286288 49608 286340
rect 49660 286328 49666 286340
rect 180702 286328 180708 286340
rect 49660 286300 180708 286328
rect 49660 286288 49666 286300
rect 180702 286288 180708 286300
rect 180760 286288 180766 286340
rect 133782 286220 133788 286272
rect 133840 286260 133846 286272
rect 186682 286260 186688 286272
rect 133840 286232 186688 286260
rect 133840 286220 133846 286232
rect 186682 286220 186688 286232
rect 186740 286220 186746 286272
rect 132310 286152 132316 286204
rect 132368 286192 132374 286204
rect 186774 286192 186780 286204
rect 132368 286164 186780 286192
rect 132368 286152 132374 286164
rect 186774 286152 186780 286164
rect 186832 286152 186838 286204
rect 126882 286084 126888 286136
rect 126940 286124 126946 286136
rect 186958 286124 186964 286136
rect 126940 286096 186964 286124
rect 126940 286084 126946 286096
rect 186958 286084 186964 286096
rect 187016 286084 187022 286136
rect 111702 286016 111708 286068
rect 111760 286056 111766 286068
rect 191374 286056 191380 286068
rect 111760 286028 191380 286056
rect 111760 286016 111766 286028
rect 191374 286016 191380 286028
rect 191432 286016 191438 286068
rect 108942 285948 108948 286000
rect 109000 285988 109006 286000
rect 188798 285988 188804 286000
rect 109000 285960 188804 285988
rect 109000 285948 109006 285960
rect 188798 285948 188804 285960
rect 188856 285948 188862 286000
rect 104802 285880 104808 285932
rect 104860 285920 104866 285932
rect 187326 285920 187332 285932
rect 104860 285892 187332 285920
rect 104860 285880 104866 285892
rect 187326 285880 187332 285892
rect 187384 285880 187390 285932
rect 86862 285812 86868 285864
rect 86920 285852 86926 285864
rect 188338 285852 188344 285864
rect 86920 285824 188344 285852
rect 86920 285812 86926 285824
rect 188338 285812 188344 285824
rect 188396 285812 188402 285864
rect 81342 285744 81348 285796
rect 81400 285784 81406 285796
rect 196710 285784 196716 285796
rect 81400 285756 196716 285784
rect 81400 285744 81406 285756
rect 196710 285744 196716 285756
rect 196768 285744 196774 285796
rect 79962 285676 79968 285728
rect 80020 285716 80026 285728
rect 196618 285716 196624 285728
rect 80020 285688 196624 285716
rect 80020 285676 80026 285688
rect 196618 285676 196624 285688
rect 196676 285676 196682 285728
rect 234982 285676 234988 285728
rect 235040 285716 235046 285728
rect 237466 285716 237472 285728
rect 235040 285688 237472 285716
rect 235040 285676 235046 285688
rect 237466 285676 237472 285688
rect 237524 285676 237530 285728
rect 113818 285608 113824 285660
rect 113876 285648 113882 285660
rect 188890 285648 188896 285660
rect 113876 285620 188896 285648
rect 113876 285608 113882 285620
rect 188890 285608 188896 285620
rect 188948 285608 188954 285660
rect 106182 285540 106188 285592
rect 106240 285580 106246 285592
rect 188706 285580 188712 285592
rect 106240 285552 188712 285580
rect 106240 285540 106246 285552
rect 188706 285540 188712 285552
rect 188764 285540 188770 285592
rect 102042 285472 102048 285524
rect 102100 285512 102106 285524
rect 195238 285512 195244 285524
rect 102100 285484 195244 285512
rect 102100 285472 102106 285484
rect 195238 285472 195244 285484
rect 195296 285472 195302 285524
rect 96154 285404 96160 285456
rect 96212 285444 96218 285456
rect 193950 285444 193956 285456
rect 96212 285416 193956 285444
rect 96212 285404 96218 285416
rect 193950 285404 193956 285416
rect 194008 285404 194014 285456
rect 93670 285336 93676 285388
rect 93728 285376 93734 285388
rect 191282 285376 191288 285388
rect 93728 285348 191288 285376
rect 93728 285336 93734 285348
rect 191282 285336 191288 285348
rect 191340 285336 191346 285388
rect 89622 285268 89628 285320
rect 89680 285308 89686 285320
rect 189902 285308 189908 285320
rect 89680 285280 189908 285308
rect 89680 285268 89686 285280
rect 189902 285268 189908 285280
rect 189960 285268 189966 285320
rect 128722 285200 128728 285252
rect 128780 285240 128786 285252
rect 238662 285240 238668 285252
rect 128780 285212 238668 285240
rect 128780 285200 128786 285212
rect 238662 285200 238668 285212
rect 238720 285200 238726 285252
rect 123570 285132 123576 285184
rect 123628 285172 123634 285184
rect 238110 285172 238116 285184
rect 123628 285144 238116 285172
rect 123628 285132 123634 285144
rect 238110 285132 238116 285144
rect 238168 285132 238174 285184
rect 118602 285064 118608 285116
rect 118660 285104 118666 285116
rect 238386 285104 238392 285116
rect 118660 285076 238392 285104
rect 118660 285064 118666 285076
rect 238386 285064 238392 285076
rect 238444 285064 238450 285116
rect 98546 284996 98552 285048
rect 98604 285036 98610 285048
rect 238478 285036 238484 285048
rect 98604 285008 238484 285036
rect 98604 284996 98610 285008
rect 238478 284996 238484 285008
rect 238536 284996 238542 285048
rect 91186 284928 91192 284980
rect 91244 284968 91250 284980
rect 238018 284968 238024 284980
rect 91244 284940 238024 284968
rect 91244 284928 91250 284940
rect 238018 284928 238024 284940
rect 238076 284928 238082 284980
rect 169754 284860 169760 284912
rect 169812 284900 169818 284912
rect 238202 284900 238208 284912
rect 169812 284872 238208 284900
rect 169812 284860 169818 284872
rect 238202 284860 238208 284872
rect 238260 284860 238266 284912
rect 232866 284316 232872 284368
rect 232924 284356 232930 284368
rect 237374 284356 237380 284368
rect 232924 284328 237380 284356
rect 232924 284316 232930 284328
rect 237374 284316 237380 284328
rect 237432 284316 237438 284368
rect 137278 283568 137284 283620
rect 137336 283608 137342 283620
rect 238570 283608 238576 283620
rect 137336 283580 238576 283608
rect 137336 283568 137342 283580
rect 238570 283568 238576 283580
rect 238628 283568 238634 283620
rect 232774 282888 232780 282940
rect 232832 282928 232838 282940
rect 237466 282928 237472 282940
rect 232832 282900 237472 282928
rect 232832 282888 232838 282900
rect 237466 282888 237472 282900
rect 237524 282888 237530 282940
rect 186682 282820 186688 282872
rect 186740 282860 186746 282872
rect 237374 282860 237380 282872
rect 186740 282832 237380 282860
rect 186740 282820 186746 282832
rect 237374 282820 237380 282832
rect 237432 282820 237438 282872
rect 196802 281528 196808 281580
rect 196860 281568 196866 281580
rect 237374 281568 237380 281580
rect 196860 281540 237380 281568
rect 196860 281528 196866 281540
rect 237374 281528 237380 281540
rect 237432 281528 237438 281580
rect 191190 280168 191196 280220
rect 191248 280208 191254 280220
rect 237466 280208 237472 280220
rect 191248 280180 237472 280208
rect 191248 280168 191254 280180
rect 237466 280168 237472 280180
rect 237524 280168 237530 280220
rect 186774 280100 186780 280152
rect 186832 280140 186838 280152
rect 237374 280140 237380 280152
rect 186832 280112 237380 280140
rect 186832 280100 186838 280112
rect 237374 280100 237380 280112
rect 237432 280100 237438 280152
rect 189074 278740 189080 278792
rect 189132 278780 189138 278792
rect 192570 278780 192576 278792
rect 189132 278752 192576 278780
rect 189132 278740 189138 278752
rect 192570 278740 192576 278752
rect 192628 278740 192634 278792
rect 189810 274728 189816 274780
rect 189868 274768 189874 274780
rect 237374 274768 237380 274780
rect 189868 274740 237380 274768
rect 189868 274728 189874 274740
rect 237374 274728 237380 274740
rect 237432 274728 237438 274780
rect 188430 274660 188436 274712
rect 188488 274700 188494 274712
rect 237466 274700 237472 274712
rect 188488 274672 237472 274700
rect 188488 274660 188494 274672
rect 237466 274660 237472 274672
rect 237524 274660 237530 274712
rect 186958 274592 186964 274644
rect 187016 274632 187022 274644
rect 237374 274632 237380 274644
rect 187016 274604 237380 274632
rect 187016 274592 187022 274604
rect 237374 274592 237380 274604
rect 237432 274592 237438 274644
rect 186958 271872 186964 271924
rect 187016 271912 187022 271924
rect 237374 271912 237380 271924
rect 187016 271884 237380 271912
rect 187016 271872 187022 271884
rect 237374 271872 237380 271884
rect 237432 271872 237438 271924
rect 540330 271872 540336 271924
rect 540388 271912 540394 271924
rect 580166 271912 580172 271924
rect 540388 271884 580172 271912
rect 540388 271872 540394 271884
rect 580166 271872 580172 271884
rect 580224 271872 580230 271924
rect 188522 269084 188528 269136
rect 188580 269124 188586 269136
rect 237374 269124 237380 269136
rect 188580 269096 237380 269124
rect 188580 269084 188586 269096
rect 237374 269084 237380 269096
rect 237432 269084 237438 269136
rect 189994 264936 190000 264988
rect 190052 264976 190058 264988
rect 237374 264976 237380 264988
rect 190052 264948 237380 264976
rect 190052 264936 190058 264948
rect 237374 264936 237380 264948
rect 237432 264936 237438 264988
rect 188614 262216 188620 262268
rect 188672 262256 188678 262268
rect 237374 262256 237380 262268
rect 188672 262228 237380 262256
rect 188672 262216 188678 262228
rect 237374 262216 237380 262228
rect 237432 262216 237438 262268
rect 193858 259496 193864 259548
rect 193916 259536 193922 259548
rect 237374 259536 237380 259548
rect 193916 259508 237380 259536
rect 193916 259496 193922 259508
rect 237374 259496 237380 259508
rect 237432 259496 237438 259548
rect 187050 259428 187056 259480
rect 187108 259468 187114 259480
rect 237466 259468 237472 259480
rect 187108 259440 237472 259468
rect 187108 259428 187114 259440
rect 237466 259428 237472 259440
rect 237524 259428 237530 259480
rect 188890 259360 188896 259412
rect 188948 259400 188954 259412
rect 237374 259400 237380 259412
rect 188948 259372 237380 259400
rect 188948 259360 188954 259372
rect 237374 259360 237380 259372
rect 237432 259360 237438 259412
rect 191374 256640 191380 256692
rect 191432 256680 191438 256692
rect 237466 256680 237472 256692
rect 191432 256652 237472 256680
rect 191432 256640 191438 256652
rect 237466 256640 237472 256652
rect 237524 256640 237530 256692
rect 192754 255280 192760 255332
rect 192812 255320 192818 255332
rect 237374 255320 237380 255332
rect 192812 255292 237380 255320
rect 192812 255280 192818 255292
rect 237374 255280 237380 255292
rect 237432 255280 237438 255332
rect 187142 253920 187148 253972
rect 187200 253960 187206 253972
rect 237374 253960 237380 253972
rect 187200 253932 237380 253960
rect 187200 253920 187206 253932
rect 237374 253920 237380 253932
rect 237432 253920 237438 253972
rect 190086 252560 190092 252612
rect 190144 252600 190150 252612
rect 237466 252600 237472 252612
rect 190144 252572 237472 252600
rect 190144 252560 190150 252572
rect 237466 252560 237472 252572
rect 237524 252560 237530 252612
rect 188798 252492 188804 252544
rect 188856 252532 188862 252544
rect 237374 252532 237380 252544
rect 188856 252504 237380 252532
rect 188856 252492 188862 252504
rect 237374 252492 237380 252504
rect 237432 252492 237438 252544
rect 191374 249772 191380 249824
rect 191432 249812 191438 249824
rect 237374 249812 237380 249824
rect 191432 249784 237380 249812
rect 191432 249772 191438 249784
rect 237374 249772 237380 249784
rect 237432 249772 237438 249824
rect 188706 248344 188712 248396
rect 188764 248384 188770 248396
rect 237374 248384 237380 248396
rect 188764 248356 237380 248384
rect 188764 248344 188770 248356
rect 237374 248344 237380 248356
rect 237432 248344 237438 248396
rect 187234 245624 187240 245676
rect 187292 245664 187298 245676
rect 237374 245664 237380 245676
rect 187292 245636 237380 245664
rect 187292 245624 187298 245636
rect 237374 245624 237380 245636
rect 237432 245624 237438 245676
rect 194042 244264 194048 244316
rect 194100 244304 194106 244316
rect 237374 244304 237380 244316
rect 194100 244276 237380 244304
rect 194100 244264 194106 244276
rect 237374 244264 237380 244276
rect 237432 244264 237438 244316
rect 187326 242836 187332 242888
rect 187384 242876 187390 242888
rect 237374 242876 237380 242888
rect 187384 242848 237380 242876
rect 187384 242836 187390 242848
rect 237374 242836 237380 242848
rect 237432 242836 237438 242888
rect 3234 240116 3240 240168
rect 3292 240156 3298 240168
rect 46290 240156 46296 240168
rect 3292 240128 46296 240156
rect 3292 240116 3298 240128
rect 46290 240116 46296 240128
rect 46348 240116 46354 240168
rect 190178 240116 190184 240168
rect 190236 240156 190242 240168
rect 237374 240156 237380 240168
rect 190236 240128 237380 240156
rect 190236 240116 190242 240128
rect 237374 240116 237380 240128
rect 237432 240116 237438 240168
rect 195238 237328 195244 237380
rect 195296 237368 195302 237380
rect 237374 237368 237380 237380
rect 195296 237340 237380 237368
rect 195296 237328 195302 237340
rect 237374 237328 237380 237340
rect 237432 237328 237438 237380
rect 188706 235968 188712 236020
rect 188764 236008 188770 236020
rect 237374 236008 237380 236020
rect 188764 235980 237380 236008
rect 188764 235968 188770 235980
rect 237374 235968 237380 235980
rect 237432 235968 237438 236020
rect 540422 231820 540428 231872
rect 540480 231860 540486 231872
rect 580166 231860 580172 231872
rect 540480 231832 580172 231860
rect 540480 231820 540486 231832
rect 580166 231820 580172 231832
rect 580224 231820 580230 231872
rect 188798 230460 188804 230512
rect 188856 230500 188862 230512
rect 237374 230500 237380 230512
rect 188856 230472 237380 230500
rect 188856 230460 188862 230472
rect 237374 230460 237380 230472
rect 237432 230460 237438 230512
rect 235810 227808 235816 227860
rect 235868 227848 235874 227860
rect 237374 227848 237380 227860
rect 235868 227820 237380 227848
rect 235868 227808 235874 227820
rect 237374 227808 237380 227820
rect 237432 227808 237438 227860
rect 195238 227740 195244 227792
rect 195296 227780 195302 227792
rect 237466 227780 237472 227792
rect 195296 227752 237472 227780
rect 195296 227740 195302 227752
rect 237466 227740 237472 227752
rect 237524 227740 237530 227792
rect 193950 227672 193956 227724
rect 194008 227712 194014 227724
rect 237374 227712 237380 227724
rect 194008 227684 237380 227712
rect 194008 227672 194014 227684
rect 237374 227672 237380 227684
rect 237432 227672 237438 227724
rect 191466 224952 191472 225004
rect 191524 224992 191530 225004
rect 237374 224992 237380 225004
rect 191524 224964 237380 224992
rect 191524 224952 191530 224964
rect 237374 224952 237380 224964
rect 237432 224952 237438 225004
rect 193950 223592 193956 223644
rect 194008 223632 194014 223644
rect 237374 223632 237380 223644
rect 194008 223604 237380 223632
rect 194008 223592 194014 223604
rect 237374 223592 237380 223604
rect 237432 223592 237438 223644
rect 191282 222096 191288 222148
rect 191340 222136 191346 222148
rect 237374 222136 237380 222148
rect 191340 222108 237380 222136
rect 191340 222096 191346 222108
rect 237374 222096 237380 222108
rect 237432 222096 237438 222148
rect 188890 220804 188896 220856
rect 188948 220844 188954 220856
rect 237374 220844 237380 220856
rect 188948 220816 237380 220844
rect 188948 220804 188954 220816
rect 237374 220804 237380 220816
rect 237432 220804 237438 220856
rect 189074 218084 189080 218136
rect 189132 218124 189138 218136
rect 192846 218124 192852 218136
rect 189132 218096 192852 218124
rect 189132 218084 189138 218096
rect 192846 218084 192852 218096
rect 192904 218084 192910 218136
rect 193122 218016 193128 218068
rect 193180 218056 193186 218068
rect 237374 218056 237380 218068
rect 193180 218028 237380 218056
rect 193180 218016 193186 218028
rect 237374 218016 237380 218028
rect 237432 218016 237438 218068
rect 190270 216724 190276 216776
rect 190328 216764 190334 216776
rect 237374 216764 237380 216776
rect 190328 216736 237380 216764
rect 190328 216724 190334 216736
rect 237374 216724 237380 216736
rect 237432 216724 237438 216776
rect 189074 216656 189080 216708
rect 189132 216696 189138 216708
rect 191282 216696 191288 216708
rect 189132 216668 191288 216696
rect 189132 216656 189138 216668
rect 191282 216656 191288 216668
rect 191340 216656 191346 216708
rect 189166 215364 189172 215416
rect 189224 215404 189230 215416
rect 191558 215404 191564 215416
rect 189224 215376 191564 215404
rect 189224 215364 189230 215376
rect 191558 215364 191564 215376
rect 191616 215364 191622 215416
rect 188982 215296 188988 215348
rect 189040 215336 189046 215348
rect 237374 215336 237380 215348
rect 189040 215308 237380 215336
rect 189040 215296 189046 215308
rect 237374 215296 237380 215308
rect 237432 215296 237438 215348
rect 187326 213936 187332 213988
rect 187384 213976 187390 213988
rect 237466 213976 237472 213988
rect 187384 213948 237472 213976
rect 187384 213936 187390 213948
rect 237466 213936 237472 213948
rect 237524 213936 237530 213988
rect 190454 213868 190460 213920
rect 190512 213908 190518 213920
rect 237374 213908 237380 213920
rect 190512 213880 237380 213908
rect 190512 213868 190518 213880
rect 237374 213868 237380 213880
rect 237432 213868 237438 213920
rect 189074 213800 189080 213852
rect 189132 213840 189138 213852
rect 193122 213840 193128 213852
rect 189132 213812 193128 213840
rect 189132 213800 189138 213812
rect 193122 213800 193128 213812
rect 193180 213800 193186 213852
rect 190362 212508 190368 212560
rect 190420 212548 190426 212560
rect 237374 212548 237380 212560
rect 190420 212520 237380 212548
rect 190420 212508 190426 212520
rect 237374 212508 237380 212520
rect 237432 212508 237438 212560
rect 189902 212440 189908 212492
rect 189960 212480 189966 212492
rect 237466 212480 237472 212492
rect 189960 212452 237472 212480
rect 189960 212440 189966 212452
rect 237466 212440 237472 212452
rect 237524 212440 237530 212492
rect 188246 209856 188252 209908
rect 188304 209896 188310 209908
rect 237466 209896 237472 209908
rect 188304 209868 237472 209896
rect 188304 209856 188310 209868
rect 237466 209856 237472 209868
rect 237524 209856 237530 209908
rect 187418 209788 187424 209840
rect 187476 209828 187482 209840
rect 237374 209828 237380 209840
rect 187476 209800 237380 209828
rect 187476 209788 187482 209800
rect 237374 209788 237380 209800
rect 237432 209788 237438 209840
rect 191558 209720 191564 209772
rect 191616 209760 191622 209772
rect 237466 209760 237472 209772
rect 191616 209732 237472 209760
rect 191616 209720 191622 209732
rect 237466 209720 237472 209732
rect 237524 209720 237530 209772
rect 47578 207680 47584 207732
rect 47636 207720 47642 207732
rect 48222 207720 48228 207732
rect 47636 207692 48228 207720
rect 47636 207680 47642 207692
rect 48222 207680 48228 207692
rect 48280 207720 48286 207732
rect 49602 207720 49608 207732
rect 48280 207692 49608 207720
rect 48280 207680 48286 207692
rect 49602 207680 49608 207692
rect 49660 207680 49666 207732
rect 189626 207000 189632 207052
rect 189684 207040 189690 207052
rect 237374 207040 237380 207052
rect 189684 207012 237380 207040
rect 189684 207000 189690 207012
rect 237374 207000 237380 207012
rect 237432 207000 237438 207052
rect 188338 206932 188344 206984
rect 188396 206972 188402 206984
rect 237466 206972 237472 206984
rect 188396 206944 237472 206972
rect 188396 206932 188402 206944
rect 237466 206932 237472 206944
rect 237524 206932 237530 206984
rect 188154 205640 188160 205692
rect 188212 205680 188218 205692
rect 237374 205680 237380 205692
rect 188212 205652 237380 205680
rect 188212 205640 188218 205652
rect 237374 205640 237380 205652
rect 237432 205640 237438 205692
rect 191282 202784 191288 202836
rect 191340 202824 191346 202836
rect 237374 202824 237380 202836
rect 191340 202796 237380 202824
rect 191340 202784 191346 202796
rect 237374 202784 237380 202796
rect 237432 202784 237438 202836
rect 189074 201492 189080 201544
rect 189132 201532 189138 201544
rect 237374 201532 237380 201544
rect 189132 201504 237380 201532
rect 189132 201492 189138 201504
rect 237374 201492 237380 201504
rect 237432 201492 237438 201544
rect 186958 200744 186964 200796
rect 187016 200784 187022 200796
rect 238202 200784 238208 200796
rect 187016 200756 238208 200784
rect 187016 200744 187022 200756
rect 238202 200744 238208 200756
rect 238260 200744 238266 200796
rect 188338 200132 188344 200184
rect 188396 200172 188402 200184
rect 237374 200172 237380 200184
rect 188396 200144 237380 200172
rect 188396 200132 188402 200144
rect 237374 200132 237380 200144
rect 237432 200132 237438 200184
rect 128354 199520 128360 199572
rect 128412 199560 128418 199572
rect 238110 199560 238116 199572
rect 128412 199532 238116 199560
rect 128412 199520 128418 199532
rect 238110 199520 238116 199532
rect 238168 199520 238174 199572
rect 120074 199452 120080 199504
rect 120132 199492 120138 199504
rect 237834 199492 237840 199504
rect 120132 199464 237840 199492
rect 120132 199452 120138 199464
rect 237834 199452 237840 199464
rect 237892 199452 237898 199504
rect 110414 199384 110420 199436
rect 110472 199424 110478 199436
rect 238018 199424 238024 199436
rect 110472 199396 238024 199424
rect 110472 199384 110478 199396
rect 238018 199384 238024 199396
rect 238076 199384 238082 199436
rect 111058 199316 111064 199368
rect 111116 199356 111122 199368
rect 187142 199356 187148 199368
rect 111116 199328 187148 199356
rect 111116 199316 111122 199328
rect 187142 199316 187148 199328
rect 187200 199316 187206 199368
rect 91186 199248 91192 199300
rect 91244 199288 91250 199300
rect 188982 199288 188988 199300
rect 91244 199260 188988 199288
rect 91244 199248 91250 199260
rect 188982 199248 188988 199260
rect 189040 199248 189046 199300
rect 88610 199180 88616 199232
rect 88668 199220 88674 199232
rect 188246 199220 188252 199232
rect 88668 199192 188252 199220
rect 88668 199180 88674 199192
rect 188246 199180 188252 199192
rect 188304 199180 188310 199232
rect 78858 199112 78864 199164
rect 78916 199152 78922 199164
rect 187326 199152 187332 199164
rect 78916 199124 187332 199152
rect 78916 199112 78922 199124
rect 187326 199112 187332 199124
rect 187384 199112 187390 199164
rect 77754 199044 77760 199096
rect 77812 199084 77818 199096
rect 187418 199084 187424 199096
rect 77812 199056 187424 199084
rect 77812 199044 77818 199056
rect 187418 199044 187424 199056
rect 187476 199044 187482 199096
rect 70578 198976 70584 199028
rect 70636 199016 70642 199028
rect 188338 199016 188344 199028
rect 70636 198988 188344 199016
rect 70636 198976 70642 198988
rect 188338 198976 188344 198988
rect 188396 198976 188402 199028
rect 103698 198908 103704 198960
rect 103756 198948 103762 198960
rect 238570 198948 238576 198960
rect 103756 198920 238576 198948
rect 103756 198908 103762 198920
rect 238570 198908 238576 198920
rect 238628 198908 238634 198960
rect 82538 198840 82544 198892
rect 82596 198880 82602 198892
rect 238478 198880 238484 198892
rect 82596 198852 238484 198880
rect 82596 198840 82602 198852
rect 238478 198840 238484 198852
rect 238536 198840 238542 198892
rect 80146 198772 80152 198824
rect 80204 198812 80210 198824
rect 238294 198812 238300 198824
rect 80204 198784 238300 198812
rect 80204 198772 80210 198784
rect 238294 198772 238300 198784
rect 238352 198772 238358 198824
rect 81342 198704 81348 198756
rect 81400 198744 81406 198756
rect 238662 198744 238668 198756
rect 81400 198716 238668 198744
rect 81400 198704 81406 198716
rect 238662 198704 238668 198716
rect 238720 198704 238726 198756
rect 86218 198636 86224 198688
rect 86276 198676 86282 198688
rect 110414 198676 110420 198688
rect 86276 198648 110420 198676
rect 86276 198636 86282 198648
rect 110414 198636 110420 198648
rect 110472 198636 110478 198688
rect 120994 198636 121000 198688
rect 121052 198676 121058 198688
rect 128354 198676 128360 198688
rect 121052 198648 128360 198676
rect 121052 198636 121058 198648
rect 128354 198636 128360 198648
rect 128412 198636 128418 198688
rect 105906 198568 105912 198620
rect 105964 198608 105970 198620
rect 235626 198608 235632 198620
rect 105964 198580 235632 198608
rect 105964 198568 105970 198580
rect 235626 198568 235632 198580
rect 235684 198568 235690 198620
rect 108482 198500 108488 198552
rect 108540 198540 108546 198552
rect 238386 198540 238392 198552
rect 108540 198512 238392 198540
rect 108540 198500 108546 198512
rect 238386 198500 238392 198512
rect 238444 198500 238450 198552
rect 71866 198432 71872 198484
rect 71924 198472 71930 198484
rect 188154 198472 188160 198484
rect 71924 198444 188160 198472
rect 71924 198432 71930 198444
rect 188154 198432 188160 198444
rect 188212 198432 188218 198484
rect 92842 198364 92848 198416
rect 92900 198404 92906 198416
rect 189994 198404 190000 198416
rect 92900 198376 190000 198404
rect 92900 198364 92906 198376
rect 189994 198364 190000 198376
rect 190052 198364 190058 198416
rect 93578 198296 93584 198348
rect 93636 198336 93642 198348
rect 188890 198336 188896 198348
rect 93636 198308 188896 198336
rect 93636 198296 93642 198308
rect 188890 198296 188896 198308
rect 188948 198296 188954 198348
rect 95970 198228 95976 198280
rect 96028 198268 96034 198280
rect 191466 198268 191472 198280
rect 96028 198240 191472 198268
rect 96028 198228 96034 198240
rect 191466 198228 191472 198240
rect 191524 198228 191530 198280
rect 98362 198160 98368 198212
rect 98420 198200 98426 198212
rect 188798 198200 188804 198212
rect 98420 198172 188804 198200
rect 98420 198160 98426 198172
rect 188798 198160 188804 198172
rect 188856 198160 188862 198212
rect 100938 198092 100944 198144
rect 100996 198132 101002 198144
rect 188706 198132 188712 198144
rect 100996 198104 188712 198132
rect 100996 198092 101002 198104
rect 188706 198092 188712 198104
rect 188764 198092 188770 198144
rect 106090 198024 106096 198076
rect 106148 198064 106154 198076
rect 187234 198064 187240 198076
rect 106148 198036 187240 198064
rect 106148 198024 106154 198036
rect 187234 198024 187240 198036
rect 187292 198024 187298 198076
rect 75546 197956 75552 198008
rect 75604 197996 75610 198008
rect 237374 197996 237380 198008
rect 75604 197968 237380 197996
rect 75604 197956 75610 197968
rect 237374 197956 237380 197968
rect 237432 197956 237438 198008
rect 113634 197888 113640 197940
rect 113692 197928 113698 197940
rect 186958 197928 186964 197940
rect 113692 197900 186964 197928
rect 113692 197888 113698 197900
rect 186958 197888 186964 197900
rect 187016 197888 187022 197940
rect 76834 197820 76840 197872
rect 76892 197860 76898 197872
rect 120074 197860 120080 197872
rect 76892 197832 120080 197860
rect 76892 197820 76898 197832
rect 120074 197820 120080 197832
rect 120132 197820 120138 197872
rect 123570 197820 123576 197872
rect 123628 197860 123634 197872
rect 188522 197860 188528 197872
rect 123628 197832 188528 197860
rect 123628 197820 123634 197832
rect 188522 197820 188528 197832
rect 188580 197820 188586 197872
rect 128906 197752 128912 197804
rect 128964 197792 128970 197804
rect 188430 197792 188436 197804
rect 128964 197764 188436 197792
rect 128964 197752 128970 197764
rect 188430 197752 188436 197764
rect 188488 197752 188494 197804
rect 47946 197684 47952 197736
rect 48004 197724 48010 197736
rect 237926 197724 237932 197736
rect 48004 197696 237932 197724
rect 48004 197684 48010 197696
rect 237926 197684 237932 197696
rect 237984 197684 237990 197736
rect 173434 197276 173440 197328
rect 173492 197316 173498 197328
rect 195238 197316 195244 197328
rect 173492 197288 195244 197316
rect 173492 197276 173498 197288
rect 195238 197276 195244 197288
rect 195296 197276 195302 197328
rect 48038 197208 48044 197260
rect 48096 197248 48102 197260
rect 190270 197248 190276 197260
rect 48096 197220 190276 197248
rect 48096 197208 48102 197220
rect 190270 197208 190276 197220
rect 190328 197208 190334 197260
rect 192846 197208 192852 197260
rect 192904 197248 192910 197260
rect 237374 197248 237380 197260
rect 192904 197220 237380 197248
rect 192904 197208 192910 197220
rect 237374 197208 237380 197220
rect 237432 197208 237438 197260
rect 85850 197140 85856 197192
rect 85908 197180 85914 197192
rect 194042 197180 194048 197192
rect 85908 197152 194048 197180
rect 85908 197140 85914 197152
rect 194042 197140 194048 197152
rect 194100 197140 194106 197192
rect 84562 197072 84568 197124
rect 84620 197112 84626 197124
rect 190178 197112 190184 197124
rect 84620 197084 190184 197112
rect 84620 197072 84626 197084
rect 190178 197072 190184 197084
rect 190236 197072 190242 197124
rect 87966 197004 87972 197056
rect 88024 197044 88030 197056
rect 191374 197044 191380 197056
rect 88024 197016 191380 197044
rect 88024 197004 88030 197016
rect 191374 197004 191380 197016
rect 191432 197004 191438 197056
rect 89530 196936 89536 196988
rect 89588 196976 89594 196988
rect 192754 196976 192760 196988
rect 89588 196948 192760 196976
rect 89588 196936 89594 196948
rect 192754 196936 192760 196948
rect 192812 196936 192818 196988
rect 90818 196868 90824 196920
rect 90876 196908 90882 196920
rect 193858 196908 193864 196920
rect 90876 196880 193864 196908
rect 90876 196868 90882 196880
rect 193858 196868 193864 196880
rect 193916 196868 193922 196920
rect 88242 196800 88248 196852
rect 88300 196840 88306 196852
rect 190086 196840 190092 196852
rect 88300 196812 190092 196840
rect 88300 196800 88306 196812
rect 190086 196800 190092 196812
rect 190144 196800 190150 196852
rect 118418 196732 118424 196784
rect 118476 196772 118482 196784
rect 188614 196772 188620 196784
rect 118476 196744 188620 196772
rect 118476 196732 118482 196744
rect 188614 196732 188620 196744
rect 188672 196732 188678 196784
rect 117038 196664 117044 196716
rect 117096 196704 117102 196716
rect 187050 196704 187056 196716
rect 117096 196676 187056 196704
rect 117096 196664 117102 196676
rect 187050 196664 187056 196676
rect 187108 196664 187114 196716
rect 73430 196596 73436 196648
rect 73488 196636 73494 196648
rect 238018 196636 238024 196648
rect 73488 196608 238024 196636
rect 73488 196596 73494 196608
rect 238018 196596 238024 196608
rect 238076 196596 238082 196648
rect 126606 196528 126612 196580
rect 126664 196568 126670 196580
rect 186866 196568 186872 196580
rect 126664 196540 186872 196568
rect 126664 196528 126670 196540
rect 186866 196528 186872 196540
rect 186924 196528 186930 196580
rect 83642 196460 83648 196512
rect 83700 196500 83706 196512
rect 237466 196500 237472 196512
rect 83700 196472 237472 196500
rect 83700 196460 83706 196472
rect 237466 196460 237472 196472
rect 237524 196460 237530 196512
rect 173250 196392 173256 196444
rect 173308 196432 173314 196444
rect 193950 196432 193956 196444
rect 173308 196404 193956 196432
rect 173308 196392 173314 196404
rect 193950 196392 193956 196404
rect 194008 196392 194014 196444
rect 49510 195916 49516 195968
rect 49568 195956 49574 195968
rect 237374 195956 237380 195968
rect 49568 195928 237380 195956
rect 49568 195916 49574 195928
rect 237374 195916 237380 195928
rect 237432 195916 237438 195968
rect 69658 195848 69664 195900
rect 69716 195888 69722 195900
rect 237466 195888 237472 195900
rect 69716 195860 237472 195888
rect 69716 195848 69722 195860
rect 237466 195848 237472 195860
rect 237524 195848 237530 195900
rect 107010 195780 107016 195832
rect 107068 195820 107074 195832
rect 235534 195820 235540 195832
rect 107068 195792 235540 195820
rect 107068 195780 107074 195792
rect 235534 195780 235540 195792
rect 235592 195780 235598 195832
rect 108574 195712 108580 195764
rect 108632 195752 108638 195764
rect 235442 195752 235448 195764
rect 108632 195724 235448 195752
rect 108632 195712 108638 195724
rect 235442 195712 235448 195724
rect 235500 195712 235506 195764
rect 109218 195644 109224 195696
rect 109276 195684 109282 195696
rect 235350 195684 235356 195696
rect 109276 195656 235356 195684
rect 109276 195644 109282 195656
rect 235350 195644 235356 195656
rect 235408 195644 235414 195696
rect 138658 195576 138664 195628
rect 138716 195616 138722 195628
rect 237098 195616 237104 195628
rect 138716 195588 237104 195616
rect 138716 195576 138722 195588
rect 237098 195576 237104 195588
rect 237156 195576 237162 195628
rect 141234 195508 141240 195560
rect 141292 195548 141298 195560
rect 237006 195548 237012 195560
rect 141292 195520 237012 195548
rect 141292 195508 141298 195520
rect 237006 195508 237012 195520
rect 237064 195508 237070 195560
rect 143442 195440 143448 195492
rect 143500 195480 143506 195492
rect 236914 195480 236920 195492
rect 143500 195452 236920 195480
rect 143500 195440 143506 195452
rect 236914 195440 236920 195452
rect 236972 195440 236978 195492
rect 146018 195372 146024 195424
rect 146076 195412 146082 195424
rect 236822 195412 236828 195424
rect 146076 195384 236828 195412
rect 146076 195372 146082 195384
rect 236822 195372 236828 195384
rect 236880 195372 236886 195424
rect 148594 195304 148600 195356
rect 148652 195344 148658 195356
rect 236730 195344 236736 195356
rect 148652 195316 236736 195344
rect 148652 195304 148658 195316
rect 236730 195304 236736 195316
rect 236788 195304 236794 195356
rect 150986 195236 150992 195288
rect 151044 195276 151050 195288
rect 232682 195276 232688 195288
rect 151044 195248 232688 195276
rect 151044 195236 151050 195248
rect 232682 195236 232688 195248
rect 232740 195236 232746 195288
rect 153378 195168 153384 195220
rect 153436 195208 153442 195220
rect 232590 195208 232596 195220
rect 153436 195180 232596 195208
rect 153436 195168 153442 195180
rect 232590 195168 232596 195180
rect 232648 195168 232654 195220
rect 133506 195100 133512 195152
rect 133564 195140 133570 195152
rect 196802 195140 196808 195152
rect 133564 195112 196808 195140
rect 133564 195100 133570 195112
rect 196802 195100 196808 195112
rect 196860 195100 196866 195152
rect 155954 194488 155960 194540
rect 156012 194528 156018 194540
rect 232498 194528 232504 194540
rect 156012 194500 232504 194528
rect 156012 194488 156018 194500
rect 232498 194488 232504 194500
rect 232556 194488 232562 194540
rect 196710 194420 196716 194472
rect 196768 194460 196774 194472
rect 237374 194460 237380 194472
rect 196768 194432 237380 194460
rect 196768 194420 196774 194432
rect 237374 194420 237380 194432
rect 237432 194420 237438 194472
rect 81250 193128 81256 193180
rect 81308 193168 81314 193180
rect 237374 193168 237380 193180
rect 81308 193140 237380 193168
rect 81308 193128 81314 193140
rect 237374 193128 237380 193140
rect 237432 193128 237438 193180
rect 74350 191768 74356 191820
rect 74408 191808 74414 191820
rect 237374 191808 237380 191820
rect 74408 191780 237380 191808
rect 74408 191768 74414 191780
rect 237374 191768 237380 191780
rect 237432 191768 237438 191820
rect 192662 191700 192668 191752
rect 192720 191740 192726 191752
rect 237466 191740 237472 191752
rect 192720 191712 237472 191740
rect 192720 191700 192726 191712
rect 237466 191700 237472 191712
rect 237524 191700 237530 191752
rect 67542 190408 67548 190460
rect 67600 190448 67606 190460
rect 237374 190448 237380 190460
rect 67600 190420 237380 190448
rect 67600 190408 67606 190420
rect 237374 190408 237380 190420
rect 237432 190408 237438 190460
rect 68922 188980 68928 189032
rect 68980 189020 68986 189032
rect 238386 189020 238392 189032
rect 68980 188992 238392 189020
rect 68980 188980 68986 188992
rect 238386 188980 238392 188992
rect 238444 188980 238450 189032
rect 3326 187688 3332 187740
rect 3384 187728 3390 187740
rect 239122 187728 239128 187740
rect 3384 187700 239128 187728
rect 3384 187688 3390 187700
rect 239122 187688 239128 187700
rect 239180 187688 239186 187740
rect 78582 187620 78588 187672
rect 78640 187660 78646 187672
rect 238754 187660 238760 187672
rect 78640 187632 238760 187660
rect 78640 187620 78646 187632
rect 238754 187620 238760 187632
rect 238812 187620 238818 187672
rect 196618 187552 196624 187604
rect 196676 187592 196682 187604
rect 238386 187592 238392 187604
rect 196676 187564 238392 187592
rect 196676 187552 196682 187564
rect 238386 187552 238392 187564
rect 238444 187552 238450 187604
rect 192478 184832 192484 184884
rect 192536 184872 192542 184884
rect 238754 184872 238760 184884
rect 192536 184844 238760 184872
rect 192536 184832 192542 184844
rect 238754 184832 238760 184844
rect 238812 184832 238818 184884
rect 49326 183472 49332 183524
rect 49384 183512 49390 183524
rect 238294 183512 238300 183524
rect 49384 183484 238300 183512
rect 49384 183472 49390 183484
rect 238294 183472 238300 183484
rect 238352 183472 238358 183524
rect 66162 183404 66168 183456
rect 66220 183444 66226 183456
rect 238386 183444 238392 183456
rect 66220 183416 238392 183444
rect 66220 183404 66226 183416
rect 238386 183404 238392 183416
rect 238444 183404 238450 183456
rect 239030 182860 239036 182912
rect 239088 182900 239094 182912
rect 239674 182900 239680 182912
rect 239088 182872 239680 182900
rect 239088 182860 239094 182872
rect 239674 182860 239680 182872
rect 239732 182860 239738 182912
rect 239306 182724 239312 182776
rect 239364 182764 239370 182776
rect 239674 182764 239680 182776
rect 239364 182736 239680 182764
rect 239364 182724 239370 182736
rect 239674 182724 239680 182736
rect 239732 182724 239738 182776
rect 192570 182112 192576 182164
rect 192628 182152 192634 182164
rect 239398 182152 239404 182164
rect 192628 182124 239404 182152
rect 192628 182112 192634 182124
rect 239398 182112 239404 182124
rect 239456 182112 239462 182164
rect 49418 181432 49424 181484
rect 49476 181472 49482 181484
rect 238570 181472 238576 181484
rect 49476 181444 238576 181472
rect 49476 181432 49482 181444
rect 238570 181432 238576 181444
rect 238628 181432 238634 181484
rect 47578 181296 47584 181348
rect 47636 181336 47642 181348
rect 48222 181336 48228 181348
rect 47636 181308 48228 181336
rect 47636 181296 47642 181308
rect 48222 181296 48228 181308
rect 48280 181296 48286 181348
rect 48222 180820 48228 180872
rect 48280 180860 48286 180872
rect 87966 180860 87972 180872
rect 48280 180832 87972 180860
rect 48280 180820 48286 180832
rect 87966 180820 87972 180832
rect 88024 180820 88030 180872
rect 300210 180208 300216 180260
rect 300268 180248 300274 180260
rect 580166 180248 580172 180260
rect 300268 180220 580172 180248
rect 300268 180208 300274 180220
rect 580166 180208 580172 180220
rect 580224 180208 580230 180260
rect 300118 180140 300124 180192
rect 300176 180180 300182 180192
rect 580902 180180 580908 180192
rect 300176 180152 580908 180180
rect 300176 180140 300182 180152
rect 580902 180140 580908 180152
rect 580960 180140 580966 180192
rect 580810 180112 580816 180124
rect 306346 180084 580816 180112
rect 297910 179868 297916 179920
rect 297968 179908 297974 179920
rect 306346 179908 306374 180084
rect 580810 180072 580816 180084
rect 580868 180072 580874 180124
rect 297968 179880 306374 179908
rect 297968 179868 297974 179880
rect 390186 179664 390192 179716
rect 390244 179704 390250 179716
rect 538306 179704 538312 179716
rect 390244 179676 538312 179704
rect 390244 179664 390250 179676
rect 538306 179664 538312 179676
rect 538364 179664 538370 179716
rect 318242 179596 318248 179648
rect 318300 179636 318306 179648
rect 540238 179636 540244 179648
rect 318300 179608 540244 179636
rect 318300 179596 318306 179608
rect 540238 179596 540244 179608
rect 540296 179596 540302 179648
rect 310330 179528 310336 179580
rect 310388 179568 310394 179580
rect 540330 179568 540336 179580
rect 310388 179540 540336 179568
rect 310388 179528 310394 179540
rect 540330 179528 540336 179540
rect 540388 179528 540394 179580
rect 302234 179460 302240 179512
rect 302292 179500 302298 179512
rect 540422 179500 540428 179512
rect 302292 179472 540428 179500
rect 302292 179460 302298 179472
rect 540422 179460 540428 179472
rect 540480 179460 540486 179512
rect 338022 179392 338028 179444
rect 338080 179432 338086 179444
rect 577498 179432 577504 179444
rect 338080 179404 577504 179432
rect 338080 179392 338086 179404
rect 577498 179392 577504 179404
rect 577556 179392 577562 179444
rect 46290 179324 46296 179376
rect 46348 179364 46354 179376
rect 517606 179364 517612 179376
rect 46348 179336 517612 179364
rect 46348 179324 46354 179336
rect 517606 179324 517612 179336
rect 517664 179324 517670 179376
rect 44818 179256 44824 179308
rect 44876 179296 44882 179308
rect 493594 179296 493600 179308
rect 44876 179268 493600 179296
rect 44876 179256 44882 179268
rect 493594 179256 493600 179268
rect 493652 179256 493658 179308
rect 46198 179188 46204 179240
rect 46256 179228 46262 179240
rect 485774 179228 485780 179240
rect 46256 179200 485780 179228
rect 46256 179188 46262 179200
rect 485774 179188 485780 179200
rect 485832 179188 485838 179240
rect 239122 179120 239128 179172
rect 239180 179160 239186 179172
rect 521654 179160 521660 179172
rect 239180 179132 521660 179160
rect 239180 179120 239186 179132
rect 521654 179120 521660 179132
rect 521712 179120 521718 179172
rect 236638 179052 236644 179104
rect 236696 179092 236702 179104
rect 509602 179092 509608 179104
rect 236696 179064 509608 179092
rect 236696 179052 236702 179064
rect 509602 179052 509608 179064
rect 509660 179052 509666 179104
rect 536926 179052 536932 179104
rect 536984 179092 536990 179104
rect 538398 179092 538404 179104
rect 536984 179064 538404 179092
rect 536984 179052 536990 179064
rect 538398 179052 538404 179064
rect 538456 179052 538462 179104
rect 233878 178984 233884 179036
rect 233936 179024 233942 179036
rect 501598 179024 501604 179036
rect 233936 178996 501604 179024
rect 233936 178984 233942 178996
rect 501598 178984 501604 178996
rect 501656 178984 501662 179036
rect 191098 178916 191104 178968
rect 191156 178956 191162 178968
rect 449986 178956 449992 178968
rect 191156 178928 449992 178956
rect 191156 178916 191162 178928
rect 449986 178916 449992 178928
rect 450044 178916 450050 178968
rect 239490 178848 239496 178900
rect 239548 178888 239554 178900
rect 477586 178888 477592 178900
rect 239548 178860 477592 178888
rect 239548 178848 239554 178860
rect 477586 178848 477592 178860
rect 477644 178848 477650 178900
rect 239858 178780 239864 178832
rect 239916 178820 239922 178832
rect 280062 178820 280068 178832
rect 239916 178792 280068 178820
rect 239916 178780 239922 178792
rect 280062 178780 280068 178792
rect 280120 178780 280126 178832
rect 355686 178780 355692 178832
rect 355744 178820 355750 178832
rect 580718 178820 580724 178832
rect 355744 178792 580724 178820
rect 355744 178780 355750 178792
rect 580718 178780 580724 178792
rect 580776 178780 580782 178832
rect 239214 178712 239220 178764
rect 239272 178752 239278 178764
rect 282914 178752 282920 178764
rect 239272 178724 282920 178752
rect 239272 178712 239278 178724
rect 282914 178712 282920 178724
rect 282972 178712 282978 178764
rect 310422 178712 310428 178764
rect 310480 178752 310486 178764
rect 580074 178752 580080 178764
rect 310480 178724 580080 178752
rect 310480 178712 310486 178724
rect 580074 178712 580080 178724
rect 580132 178712 580138 178764
rect 3694 178644 3700 178696
rect 3752 178684 3758 178696
rect 401594 178684 401600 178696
rect 3752 178656 401600 178684
rect 3752 178644 3758 178656
rect 401594 178644 401600 178656
rect 401652 178644 401658 178696
rect 408494 178644 408500 178696
rect 408552 178684 408558 178696
rect 580626 178684 580632 178696
rect 408552 178656 580632 178684
rect 408552 178644 408558 178656
rect 580626 178644 580632 178656
rect 580684 178644 580690 178696
rect 189718 178576 189724 178628
rect 189776 178616 189782 178628
rect 410058 178616 410064 178628
rect 189776 178588 410064 178616
rect 189776 178576 189782 178588
rect 410058 178576 410064 178588
rect 410116 178576 410122 178628
rect 366266 178508 366272 178560
rect 366324 178548 366330 178560
rect 580258 178548 580264 178560
rect 366324 178520 580264 178548
rect 366324 178508 366330 178520
rect 580258 178508 580264 178520
rect 580316 178508 580322 178560
rect 239674 178440 239680 178492
rect 239732 178480 239738 178492
rect 393590 178480 393596 178492
rect 239732 178452 393596 178480
rect 239732 178440 239738 178452
rect 393590 178440 393596 178452
rect 393648 178440 393654 178492
rect 406194 178032 406200 178084
rect 406252 178072 406258 178084
rect 580166 178072 580172 178084
rect 406252 178044 580172 178072
rect 406252 178032 406258 178044
rect 580166 178032 580172 178044
rect 580224 178032 580230 178084
rect 334250 177964 334256 178016
rect 334308 178004 334314 178016
rect 355686 178004 355692 178016
rect 334308 177976 355692 178004
rect 334308 177964 334314 177976
rect 355686 177964 355692 177976
rect 355744 177964 355750 178016
rect 531958 177964 531964 178016
rect 532016 178004 532022 178016
rect 538030 178004 538036 178016
rect 532016 177976 538036 178004
rect 532016 177964 532022 177976
rect 538030 177964 538036 177976
rect 538088 177964 538094 178016
rect 289906 177896 289912 177948
rect 289964 177936 289970 177948
rect 300118 177936 300124 177948
rect 289964 177908 300124 177936
rect 289964 177896 289970 177908
rect 300118 177896 300124 177908
rect 300176 177896 300182 177948
rect 3878 177828 3884 177880
rect 3936 177868 3942 177880
rect 490006 177868 490012 177880
rect 3936 177840 490012 177868
rect 3936 177828 3942 177840
rect 490006 177828 490012 177840
rect 490064 177828 490070 177880
rect 3786 177760 3792 177812
rect 3844 177800 3850 177812
rect 481634 177800 481640 177812
rect 3844 177772 481640 177800
rect 3844 177760 3850 177772
rect 481634 177760 481640 177772
rect 481692 177760 481698 177812
rect 490558 177760 490564 177812
rect 490616 177800 490622 177812
rect 513558 177800 513564 177812
rect 490616 177772 513564 177800
rect 490616 177760 490622 177772
rect 513558 177760 513564 177772
rect 513616 177760 513622 177812
rect 530670 177760 530676 177812
rect 530728 177800 530734 177812
rect 536926 177800 536932 177812
rect 530728 177772 536932 177800
rect 530728 177760 530734 177772
rect 536926 177760 536932 177772
rect 536984 177760 536990 177812
rect 87966 177692 87972 177744
rect 88024 177732 88030 177744
rect 241974 177732 241980 177744
rect 88024 177704 241980 177732
rect 88024 177692 88030 177704
rect 241974 177692 241980 177704
rect 242032 177692 242038 177744
rect 281902 177692 281908 177744
rect 281960 177732 281966 177744
rect 300210 177732 300216 177744
rect 281960 177704 300216 177732
rect 281960 177692 281966 177704
rect 300210 177692 300216 177704
rect 300268 177692 300274 177744
rect 342162 177692 342168 177744
rect 342220 177732 342226 177744
rect 580534 177732 580540 177744
rect 342220 177704 580540 177732
rect 342220 177692 342226 177704
rect 580534 177692 580540 177704
rect 580592 177692 580598 177744
rect 306190 177624 306196 177676
rect 306248 177664 306254 177676
rect 538950 177664 538956 177676
rect 306248 177636 538956 177664
rect 306248 177624 306254 177636
rect 538950 177624 538956 177636
rect 539008 177624 539014 177676
rect 293954 177556 293960 177608
rect 294012 177596 294018 177608
rect 310422 177596 310428 177608
rect 294012 177568 310428 177596
rect 294012 177556 294018 177568
rect 310422 177556 310428 177568
rect 310480 177556 310486 177608
rect 350258 177556 350264 177608
rect 350316 177596 350322 177608
rect 580442 177596 580448 177608
rect 350316 177568 580448 177596
rect 350316 177556 350322 177568
rect 580442 177556 580448 177568
rect 580500 177556 580506 177608
rect 314194 177488 314200 177540
rect 314252 177528 314258 177540
rect 538858 177528 538864 177540
rect 314252 177500 538864 177528
rect 314252 177488 314258 177500
rect 538858 177488 538864 177500
rect 538916 177488 538922 177540
rect 358170 177420 358176 177472
rect 358228 177460 358234 177472
rect 580350 177460 580356 177472
rect 358228 177432 580356 177460
rect 358228 177420 358234 177432
rect 580350 177420 580356 177432
rect 580408 177420 580414 177472
rect 362218 177352 362224 177404
rect 362276 177392 362282 177404
rect 542354 177392 542360 177404
rect 362276 177364 542360 177392
rect 362276 177352 362282 177364
rect 542354 177352 542360 177364
rect 542412 177352 542418 177404
rect 1394 177284 1400 177336
rect 1452 177324 1458 177336
rect 245930 177324 245936 177336
rect 1452 177296 245936 177324
rect 1452 177284 1458 177296
rect 245930 177284 245936 177296
rect 245988 177284 245994 177336
rect 382182 177284 382188 177336
rect 382240 177324 382246 177336
rect 538214 177324 538220 177336
rect 382240 177296 538220 177324
rect 382240 177284 382246 177296
rect 538214 177284 538220 177296
rect 538272 177284 538278 177336
rect 239030 177216 239036 177268
rect 239088 177256 239094 177268
rect 413554 177256 413560 177268
rect 239088 177228 413560 177256
rect 239088 177216 239094 177228
rect 413554 177216 413560 177228
rect 413612 177216 413618 177268
rect 273898 177148 273904 177200
rect 273956 177188 273962 177200
rect 406194 177188 406200 177200
rect 273956 177160 406200 177188
rect 273956 177148 273962 177160
rect 406194 177148 406200 177160
rect 406252 177148 406258 177200
rect 322290 177080 322296 177132
rect 322348 177120 322354 177132
rect 408494 177120 408500 177132
rect 322348 177092 408500 177120
rect 322348 177080 322354 177092
rect 408494 177080 408500 177092
rect 408552 177080 408558 177132
rect 4062 177012 4068 177064
rect 4120 177052 4126 177064
rect 505554 177052 505560 177064
rect 4120 177024 505560 177052
rect 4120 177012 4126 177024
rect 505554 177012 505560 177024
rect 505612 177012 505618 177064
rect 3970 176944 3976 176996
rect 4028 176984 4034 176996
rect 497550 176984 497556 176996
rect 4028 176956 497556 176984
rect 4028 176944 4034 176956
rect 497550 176944 497556 176956
rect 497608 176944 497614 176996
rect 3510 176604 3516 176656
rect 3568 176644 3574 176656
rect 461578 176644 461584 176656
rect 3568 176616 461584 176644
rect 3568 176604 3574 176616
rect 461578 176604 461584 176616
rect 461636 176604 461642 176656
rect 23474 176536 23480 176588
rect 23532 176576 23538 176588
rect 425606 176576 425612 176588
rect 23532 176548 425612 176576
rect 23532 176536 23538 176548
rect 425606 176536 425612 176548
rect 425664 176536 425670 176588
rect 330202 176468 330208 176520
rect 330260 176508 330266 176520
rect 577590 176508 577596 176520
rect 330260 176480 577596 176508
rect 330260 176468 330266 176480
rect 577590 176468 577596 176480
rect 577648 176468 577654 176520
rect 326338 176400 326344 176452
rect 326396 176440 326402 176452
rect 542998 176440 543004 176452
rect 326396 176412 543004 176440
rect 326396 176400 326402 176412
rect 542998 176400 543004 176412
rect 543056 176400 543062 176452
rect 378042 176332 378048 176384
rect 378100 176372 378106 176384
rect 531958 176372 531964 176384
rect 378100 176344 531964 176372
rect 378100 176332 378106 176344
rect 531958 176332 531964 176344
rect 532016 176332 532022 176384
rect 282914 176264 282920 176316
rect 282972 176304 282978 176316
rect 385586 176304 385592 176316
rect 282972 176276 385592 176304
rect 282972 176264 282978 176276
rect 385586 176264 385592 176276
rect 385644 176264 385650 176316
rect 398282 176264 398288 176316
rect 398340 176304 398346 176316
rect 530670 176304 530676 176316
rect 398340 176276 530676 176304
rect 398340 176264 398346 176276
rect 530670 176264 530676 176276
rect 530728 176264 530734 176316
rect 280062 176196 280068 176248
rect 280120 176236 280126 176248
rect 405734 176236 405740 176248
rect 280120 176208 405740 176236
rect 280120 176196 280126 176208
rect 405734 176196 405740 176208
rect 405792 176196 405798 176248
rect 235258 175176 235264 175228
rect 235316 175216 235322 175228
rect 457530 175216 457536 175228
rect 235316 175188 457536 175216
rect 235316 175176 235322 175188
rect 457530 175176 457536 175188
rect 457588 175176 457594 175228
rect 256694 174088 256700 174140
rect 256752 174128 256758 174140
rect 257890 174128 257896 174140
rect 256752 174100 257896 174128
rect 256752 174088 256758 174100
rect 257890 174088 257896 174100
rect 257948 174088 257954 174140
rect 285674 153144 285680 153196
rect 285732 153184 285738 153196
rect 580166 153184 580172 153196
rect 285732 153156 580172 153184
rect 285732 153144 285738 153156
rect 580166 153144 580172 153156
rect 580224 153144 580230 153196
rect 3418 150356 3424 150408
rect 3476 150396 3482 150408
rect 490558 150396 490564 150408
rect 3476 150368 490564 150396
rect 3476 150356 3482 150368
rect 490558 150356 490564 150368
rect 490616 150356 490622 150408
rect 264974 139340 264980 139392
rect 265032 139380 265038 139392
rect 580166 139380 580172 139392
rect 265032 139352 580172 139380
rect 265032 139340 265038 139352
rect 580166 139340 580172 139352
rect 580224 139340 580230 139392
rect 3234 137912 3240 137964
rect 3292 137952 3298 137964
rect 525794 137952 525800 137964
rect 3292 137924 525800 137952
rect 3292 137912 3298 137924
rect 525794 137912 525800 137924
rect 525852 137912 525858 137964
rect 277394 113092 277400 113144
rect 277452 113132 277458 113144
rect 579798 113132 579804 113144
rect 277452 113104 579804 113132
rect 277452 113092 277458 113104
rect 579798 113092 579804 113104
rect 579856 113092 579862 113144
rect 256694 100648 256700 100700
rect 256752 100688 256758 100700
rect 580166 100688 580172 100700
rect 256752 100660 580172 100688
rect 256752 100648 256758 100660
rect 580166 100648 580172 100660
rect 580224 100648 580230 100700
rect 3142 85484 3148 85536
rect 3200 85524 3206 85536
rect 529934 85524 529940 85536
rect 3200 85496 529940 85524
rect 3200 85484 3206 85496
rect 529934 85484 529940 85496
rect 529992 85484 529998 85536
rect 269114 73108 269120 73160
rect 269172 73148 269178 73160
rect 580166 73148 580172 73160
rect 269172 73120 580172 73148
rect 269172 73108 269178 73120
rect 580166 73108 580172 73120
rect 580224 73108 580230 73160
rect 249794 60664 249800 60716
rect 249852 60704 249858 60716
rect 580166 60704 580172 60716
rect 249852 60676 580172 60704
rect 249852 60664 249858 60676
rect 580166 60664 580172 60676
rect 580224 60664 580230 60716
rect 3418 45500 3424 45552
rect 3476 45540 3482 45552
rect 532694 45540 532700 45552
rect 3476 45512 532700 45540
rect 3476 45500 3482 45512
rect 532694 45500 532700 45512
rect 532752 45500 532758 45552
rect 260834 33056 260840 33108
rect 260892 33096 260898 33108
rect 580166 33096 580172 33108
rect 260892 33068 580172 33096
rect 260892 33056 260898 33068
rect 580166 33056 580172 33068
rect 580224 33056 580230 33108
rect 3418 6808 3424 6860
rect 3476 6848 3482 6860
rect 536834 6848 536840 6860
rect 3476 6820 536840 6848
rect 3476 6808 3482 6820
rect 536834 6808 536840 6820
rect 536892 6808 536898 6860
rect 253934 6740 253940 6792
rect 253992 6780 253998 6792
rect 580166 6780 580172 6792
rect 253992 6752 580172 6780
rect 253992 6740 253998 6752
rect 580166 6740 580172 6752
rect 580224 6740 580230 6792
rect 566 3408 572 3460
rect 624 3448 630 3460
rect 47578 3448 47584 3460
rect 624 3420 47584 3448
rect 624 3408 630 3420
rect 47578 3408 47584 3420
rect 47636 3408 47642 3460
<< via1 >>
rect 201500 702992 201552 703044
rect 202788 702992 202840 703044
rect 413652 700476 413704 700528
rect 420920 700476 420972 700528
rect 154120 700340 154172 700392
rect 189724 700340 189776 700392
rect 278780 700340 278832 700392
rect 348792 700340 348844 700392
rect 72976 700272 73028 700324
rect 239404 700272 239456 700324
rect 262220 700272 262272 700324
rect 332508 700272 332560 700324
rect 527180 700272 527232 700324
rect 538220 700272 538272 700324
rect 397460 699932 397512 699984
rect 399300 699932 399352 699984
rect 266360 697552 266412 697604
rect 267648 697552 267700 697604
rect 399300 695444 399352 695496
rect 400956 695444 401008 695496
rect 477500 694764 477552 694816
rect 480260 694764 480312 694816
rect 420920 694152 420972 694204
rect 424324 694152 424376 694204
rect 259460 694084 259512 694136
rect 262128 694084 262180 694136
rect 276756 692792 276808 692844
rect 278688 692792 278740 692844
rect 400956 691092 401008 691144
rect 401968 691092 402020 691144
rect 462320 690684 462372 690736
rect 465172 690684 465224 690736
rect 465172 688168 465224 688220
rect 471244 688168 471296 688220
rect 480260 687896 480312 687948
rect 490564 687896 490616 687948
rect 275284 687488 275336 687540
rect 276756 687488 276808 687540
rect 424324 685108 424376 685160
rect 447784 685108 447836 685160
rect 401968 684496 402020 684548
rect 405004 684428 405056 684480
rect 253204 683136 253256 683188
rect 259368 683136 259420 683188
rect 471244 681368 471296 681420
rect 474648 681368 474700 681420
rect 474648 677492 474700 677544
rect 478144 677492 478196 677544
rect 478144 672732 478196 672784
rect 483664 672732 483716 672784
rect 490564 665116 490616 665168
rect 493324 665116 493376 665168
rect 447784 664436 447836 664488
rect 460204 664436 460256 664488
rect 483664 664436 483716 664488
rect 497464 664436 497516 664488
rect 3516 656888 3568 656940
rect 239588 656888 239640 656940
rect 460204 656276 460256 656328
rect 462320 656276 462372 656328
rect 273904 655460 273956 655512
rect 275284 655460 275336 655512
rect 497464 654780 497516 654832
rect 508504 654780 508556 654832
rect 462320 653148 462372 653200
rect 465448 653148 465500 653200
rect 465448 650632 465500 650684
rect 480904 650632 480956 650684
rect 480904 641044 480956 641096
rect 494704 641044 494756 641096
rect 493324 640976 493376 641028
rect 507124 640976 507176 641028
rect 272524 638188 272576 638240
rect 273904 638188 273956 638240
rect 494704 636828 494756 636880
rect 505744 636828 505796 636880
rect 508504 633700 508556 633752
rect 511264 633700 511316 633752
rect 251824 627852 251876 627904
rect 253204 627852 253256 627904
rect 405004 626492 405056 626544
rect 407764 626492 407816 626544
rect 511264 624384 511316 624436
rect 521660 624384 521712 624436
rect 269764 623772 269816 623824
rect 272524 623772 272576 623824
rect 505744 623024 505796 623076
rect 522304 623024 522356 623076
rect 521660 616768 521712 616820
rect 525156 616768 525208 616820
rect 522304 614184 522356 614236
rect 525064 614184 525116 614236
rect 407764 613028 407816 613080
rect 409236 613028 409288 613080
rect 409236 609900 409288 609952
rect 410524 609900 410576 609952
rect 507124 607860 507176 607912
rect 518900 607860 518952 607912
rect 525156 607112 525208 607164
rect 527640 607112 527692 607164
rect 268752 604460 268804 604512
rect 269764 604460 269816 604512
rect 527640 603712 527692 603764
rect 533344 603712 533396 603764
rect 518900 603100 518952 603152
rect 522856 603100 522908 603152
rect 267004 602352 267056 602404
rect 268752 602352 268804 602404
rect 250444 600448 250496 600500
rect 251824 600448 251876 600500
rect 410524 600244 410576 600296
rect 411904 600244 411956 600296
rect 411904 595076 411956 595128
rect 414664 595076 414716 595128
rect 533344 591948 533396 592000
rect 538312 591948 538364 592000
rect 282184 588412 282236 588464
rect 282920 588412 282972 588464
rect 264980 579640 265032 579692
rect 267004 579640 267056 579692
rect 262864 578144 262916 578196
rect 264980 578144 265032 578196
rect 577504 577192 577556 577244
rect 579620 577192 579672 577244
rect 280804 575492 280856 575544
rect 282184 575492 282236 575544
rect 247684 573792 247736 573844
rect 250444 573792 250496 573844
rect 3056 565836 3108 565888
rect 191104 565836 191156 565888
rect 525064 562300 525116 562352
rect 533344 562300 533396 562352
rect 278044 561620 278096 561672
rect 280804 561688 280856 561740
rect 414664 558832 414716 558884
rect 416044 558832 416096 558884
rect 3608 553392 3660 553444
rect 239772 553392 239824 553444
rect 261208 550740 261260 550792
rect 262864 550740 262916 550792
rect 259460 548496 259512 548548
rect 261208 548496 261260 548548
rect 533344 543804 533396 543856
rect 535736 543804 535788 543856
rect 535736 542308 535788 542360
rect 538036 542308 538088 542360
rect 257344 539588 257396 539640
rect 259368 539588 259420 539640
rect 245016 532448 245068 532500
rect 247684 532448 247736 532500
rect 416044 529864 416096 529916
rect 417516 529864 417568 529916
rect 417516 526260 417568 526312
rect 418896 526260 418948 526312
rect 254584 524424 254636 524476
rect 257344 524424 257396 524476
rect 577596 524424 577648 524476
rect 579620 524424 579672 524476
rect 244924 523676 244976 523728
rect 278044 523676 278096 523728
rect 418896 521568 418948 521620
rect 420184 521568 420236 521620
rect 3332 514768 3384 514820
rect 235264 514768 235316 514820
rect 420184 514700 420236 514752
rect 422944 514700 422996 514752
rect 243636 506472 243688 506524
rect 245016 506472 245068 506524
rect 422944 505724 422996 505776
rect 424324 505724 424376 505776
rect 251640 505112 251692 505164
rect 254584 505112 254636 505164
rect 242164 504160 242216 504212
rect 243636 504160 243688 504212
rect 249800 501984 249852 502036
rect 251640 501984 251692 502036
rect 3332 500964 3384 501016
rect 239496 500964 239548 501016
rect 247684 496952 247736 497004
rect 249800 496952 249852 497004
rect 242256 496816 242308 496868
rect 244924 496816 244976 496868
rect 242808 485800 242860 485852
rect 247684 485800 247736 485852
rect 240324 484032 240376 484084
rect 242256 484032 242308 484084
rect 240784 483760 240836 483812
rect 242808 483760 242860 483812
rect 239864 482672 239916 482724
rect 242164 482672 242216 482724
rect 239680 480904 239732 480956
rect 266360 480904 266412 480956
rect 424324 480904 424376 480956
rect 437388 480904 437440 480956
rect 239220 479544 239272 479596
rect 240784 479544 240836 479596
rect 437388 479544 437440 479596
rect 538404 479476 538456 479528
rect 157248 478864 157300 478916
rect 237380 478864 237432 478916
rect 239312 478864 239364 478916
rect 240324 478864 240376 478916
rect 235540 477504 235592 477556
rect 237380 477504 237432 477556
rect 235632 476076 235684 476128
rect 237380 476076 237432 476128
rect 154488 473356 154540 473408
rect 237380 473356 237432 473408
rect 235724 472064 235776 472116
rect 237472 472064 237524 472116
rect 235816 471996 235868 472048
rect 237380 471996 237432 472048
rect 151360 469208 151412 469260
rect 237380 469208 237432 469260
rect 235908 467848 235960 467900
rect 237380 467848 237432 467900
rect 235172 466420 235224 466472
rect 237380 466420 237432 466472
rect 169760 465944 169812 465996
rect 192484 465944 192536 465996
rect 168472 465876 168524 465928
rect 192576 465876 192628 465928
rect 146024 465808 146076 465860
rect 186688 465808 186740 465860
rect 141056 465740 141108 465792
rect 187240 465740 187292 465792
rect 136088 465672 136140 465724
rect 187148 465672 187200 465724
rect 128728 465604 128780 465656
rect 187056 465604 187108 465656
rect 111064 465536 111116 465588
rect 186964 465536 187016 465588
rect 108488 465468 108540 465520
rect 188344 465468 188396 465520
rect 101312 465400 101364 465452
rect 191288 465400 191340 465452
rect 106188 465332 106240 465384
rect 198188 465332 198240 465384
rect 103704 465264 103756 465316
rect 198096 465264 198148 465316
rect 96160 465196 96212 465248
rect 191196 465196 191248 465248
rect 93676 465128 93728 465180
rect 198004 465128 198056 465180
rect 91192 465060 91244 465112
rect 235448 465060 235500 465112
rect 148508 464992 148560 465044
rect 237380 464992 237432 465044
rect 121000 464924 121052 464976
rect 189908 464924 189960 464976
rect 143632 464856 143684 464908
rect 238024 464856 238076 464908
rect 98552 464788 98604 464840
rect 199384 464788 199436 464840
rect 133512 464720 133564 464772
rect 237932 464720 237984 464772
rect 131120 464652 131172 464704
rect 238668 464652 238720 464704
rect 88524 464584 88576 464636
rect 196624 464584 196676 464636
rect 83464 464516 83516 464568
rect 193864 464516 193916 464568
rect 118608 464448 118660 464500
rect 238392 464448 238444 464500
rect 116124 464380 116176 464432
rect 238208 464380 238260 464432
rect 113640 464312 113692 464364
rect 238116 464312 238168 464364
rect 123576 464244 123628 464296
rect 190092 464244 190144 464296
rect 125968 464176 126020 464228
rect 192668 464176 192720 464228
rect 138480 464108 138532 464160
rect 188620 464108 188672 464160
rect 186688 462952 186740 463004
rect 237472 462952 237524 463004
rect 215944 462340 215996 462392
rect 237380 462340 237432 462392
rect 189080 458260 189132 458312
rect 195244 458260 195296 458312
rect 188436 458192 188488 458244
rect 237380 458192 237432 458244
rect 187240 449828 187292 449880
rect 237380 449828 237432 449880
rect 3332 448536 3384 448588
rect 46204 448536 46256 448588
rect 188528 447108 188580 447160
rect 237380 447108 237432 447160
rect 188620 444320 188672 444372
rect 237380 444320 237432 444372
rect 188620 441600 188672 441652
rect 237380 441600 237432 441652
rect 187148 440172 187200 440224
rect 237380 440172 237432 440224
rect 188712 437452 188764 437504
rect 237380 437452 237432 437504
rect 188804 431944 188856 431996
rect 237380 431944 237432 431996
rect 190000 430584 190052 430636
rect 237380 430584 237432 430636
rect 193956 426504 194008 426556
rect 237380 426504 237432 426556
rect 188896 426436 188948 426488
rect 237472 426436 237524 426488
rect 187056 423580 187108 423632
rect 237380 423580 237432 423632
rect 188988 422288 189040 422340
rect 237380 422288 237432 422340
rect 192668 419432 192720 419484
rect 237380 419432 237432 419484
rect 538956 418140 539008 418192
rect 579620 418140 579672 418192
rect 187056 416780 187108 416832
rect 237380 416780 237432 416832
rect 187148 415420 187200 415472
rect 237380 415420 237432 415472
rect 190092 413924 190144 413976
rect 237380 413924 237432 413976
rect 187240 411272 187292 411324
rect 237380 411272 237432 411324
rect 189908 408416 189960 408468
rect 237380 408416 237432 408468
rect 189908 405696 189960 405748
rect 237380 405696 237432 405748
rect 187332 401616 187384 401668
rect 237380 401616 237432 401668
rect 190092 400188 190144 400240
rect 237380 400188 237432 400240
rect 189080 398828 189132 398880
rect 192668 398828 192720 398880
rect 3332 397468 3384 397520
rect 44824 397468 44876 397520
rect 189080 397468 189132 397520
rect 192760 397468 192812 397520
rect 189080 396176 189132 396228
rect 195336 396176 195388 396228
rect 190184 396108 190236 396160
rect 237380 396108 237432 396160
rect 187424 396040 187476 396092
rect 237472 396040 237524 396092
rect 189448 394680 189500 394732
rect 195428 394680 195480 394732
rect 189080 393320 189132 393372
rect 195520 393320 195572 393372
rect 187516 391960 187568 392012
rect 237380 391960 237432 392012
rect 188252 390532 188304 390584
rect 237380 390532 237432 390584
rect 186964 389104 187016 389156
rect 237380 389104 237432 389156
rect 186964 386384 187016 386436
rect 237380 386384 237432 386436
rect 187792 385024 187844 385076
rect 237380 385024 237432 385076
rect 188344 383596 188396 383648
rect 237380 383596 237432 383648
rect 187700 380876 187752 380928
rect 237380 380876 237432 380928
rect 186688 380128 186740 380180
rect 237932 380128 237984 380180
rect 48228 379516 48280 379568
rect 49884 379516 49936 379568
rect 116032 379448 116084 379500
rect 187424 379448 187476 379500
rect 113548 379380 113600 379432
rect 187516 379380 187568 379432
rect 110972 379312 111024 379364
rect 186964 379312 187016 379364
rect 150992 379244 151044 379296
rect 235908 379244 235960 379296
rect 144920 379176 144972 379228
rect 238024 379176 238076 379228
rect 89444 379108 89496 379160
rect 188252 379108 188304 379160
rect 88156 379040 88208 379092
rect 187792 379040 187844 379092
rect 90732 378972 90784 379024
rect 190184 378972 190236 379024
rect 87052 378904 87104 378956
rect 187700 378904 187752 378956
rect 135996 378836 136048 378888
rect 237472 378836 237524 378888
rect 121000 378768 121052 378820
rect 237840 378768 237892 378820
rect 118332 378700 118384 378752
rect 187332 378700 187384 378752
rect 123484 378632 123536 378684
rect 187240 378632 187292 378684
rect 130936 378564 130988 378616
rect 188896 378564 188948 378616
rect 543004 378156 543056 378208
rect 580172 378156 580224 378208
rect 91928 378020 91980 378072
rect 190092 378020 190144 378072
rect 198188 378020 198240 378072
rect 237380 378020 237432 378072
rect 92848 377952 92900 378004
rect 189908 377952 189960 378004
rect 93952 377884 94004 377936
rect 186688 377884 186740 377936
rect 95240 377816 95292 377868
rect 187148 377816 187200 377868
rect 96436 377748 96488 377800
rect 140780 377748 140832 377800
rect 148600 377748 148652 377800
rect 215944 377748 215996 377800
rect 125968 377680 126020 377732
rect 187056 377680 187108 377732
rect 128544 377612 128596 377664
rect 188988 377612 189040 377664
rect 133512 377544 133564 377596
rect 188804 377544 188856 377596
rect 108488 377476 108540 377528
rect 135996 377476 136048 377528
rect 136088 377476 136140 377528
rect 188712 377476 188764 377528
rect 106096 377408 106148 377460
rect 237380 377408 237432 377460
rect 138664 377340 138716 377392
rect 188620 377340 188672 377392
rect 141148 377272 141200 377324
rect 188528 377272 188580 377324
rect 146024 377204 146076 377256
rect 188436 377204 188488 377256
rect 99932 377136 99984 377188
rect 238576 377136 238628 377188
rect 78312 377000 78364 377052
rect 79324 377000 79376 377052
rect 85948 376660 86000 376712
rect 237380 376660 237432 376712
rect 97632 376592 97684 376644
rect 193956 376592 194008 376644
rect 153384 376524 153436 376576
rect 235724 376524 235776 376576
rect 155960 376456 156012 376508
rect 235540 376456 235592 376508
rect 49332 375980 49384 376032
rect 238024 375980 238076 376032
rect 198096 373940 198148 373992
rect 237380 373940 237432 373992
rect 104808 372512 104860 372564
rect 237380 372512 237432 372564
rect 47860 371832 47912 371884
rect 122104 371832 122156 371884
rect 85488 371152 85540 371204
rect 237380 371152 237432 371204
rect 47952 369112 48004 369164
rect 177304 369112 177356 369164
rect 191288 368432 191340 368484
rect 237380 368432 237432 368484
rect 84016 367004 84068 367056
rect 237472 367004 237524 367056
rect 102048 366936 102100 366988
rect 237380 366936 237432 366988
rect 49424 364964 49476 365016
rect 238116 364964 238168 365016
rect 538956 364352 539008 364404
rect 580172 364352 580224 364404
rect 99288 362856 99340 362908
rect 237472 362856 237524 362908
rect 199384 362788 199436 362840
rect 237380 362788 237432 362840
rect 82728 361496 82780 361548
rect 237380 361496 237432 361548
rect 173716 360136 173768 360188
rect 237380 360136 237432 360188
rect 48044 358708 48096 358760
rect 237380 358708 237432 358760
rect 191196 358640 191248 358692
rect 237472 358640 237524 358692
rect 96528 357348 96580 357400
rect 237380 357348 237432 357400
rect 81164 355988 81216 356040
rect 237380 355988 237432 356040
rect 173808 355920 173860 355972
rect 237472 355920 237524 355972
rect 177304 354628 177356 354680
rect 237380 354628 237432 354680
rect 198004 353200 198056 353252
rect 237380 353200 237432 353252
rect 81256 351840 81308 351892
rect 237472 351840 237524 351892
rect 93768 351772 93820 351824
rect 237380 351772 237432 351824
rect 195520 350480 195572 350532
rect 237380 350480 237432 350532
rect 49884 349052 49936 349104
rect 237380 349052 237432 349104
rect 92388 347692 92440 347744
rect 237380 347692 237432 347744
rect 235448 347624 235500 347676
rect 237472 347624 237524 347676
rect 79968 346332 80020 346384
rect 237380 346332 237432 346384
rect 3056 345040 3108 345092
rect 233884 345040 233936 345092
rect 195428 344972 195480 345024
rect 237380 344972 237432 345024
rect 196624 343544 196676 343596
rect 237380 343544 237432 343596
rect 89628 342184 89680 342236
rect 237380 342184 237432 342236
rect 78496 340824 78548 340876
rect 237380 340824 237432 340876
rect 195336 340756 195388 340808
rect 237472 340756 237524 340808
rect 73068 338036 73120 338088
rect 237380 338036 237432 338088
rect 86776 336676 86828 336728
rect 237472 336676 237524 336728
rect 189816 336608 189868 336660
rect 237380 336608 237432 336660
rect 77208 335248 77260 335300
rect 237380 335248 237432 335300
rect 192760 333888 192812 333940
rect 237380 333888 237432 333940
rect 49240 332528 49292 332580
rect 237380 332528 237432 332580
rect 71688 332460 71740 332512
rect 237472 332460 237524 332512
rect 193864 331168 193916 331220
rect 237380 331168 237432 331220
rect 75828 329740 75880 329792
rect 237472 329740 237524 329792
rect 84108 329672 84160 329724
rect 237380 329672 237432 329724
rect 192668 328380 192720 328432
rect 237380 328380 237432 328432
rect 49608 327020 49660 327072
rect 237380 327020 237432 327072
rect 70308 325592 70360 325644
rect 237380 325592 237432 325644
rect 235356 325320 235408 325372
rect 237380 325320 237432 325372
rect 74356 324912 74408 324964
rect 237472 324912 237524 324964
rect 540244 324300 540296 324352
rect 579620 324300 579672 324352
rect 81348 324232 81400 324284
rect 237380 324232 237432 324284
rect 74448 323552 74500 323604
rect 237564 323552 237616 323604
rect 67548 321512 67600 321564
rect 237472 321512 237524 321564
rect 192576 321444 192628 321496
rect 237380 321444 237432 321496
rect 68928 320084 68980 320136
rect 237380 320084 237432 320136
rect 79324 317364 79376 317416
rect 237380 317364 237432 317416
rect 192484 315936 192536 315988
rect 237380 315936 237432 315988
rect 66168 314576 66220 314628
rect 237380 314576 237432 314628
rect 48136 313216 48188 313268
rect 237380 313216 237432 313268
rect 195244 313148 195296 313200
rect 237472 313148 237524 313200
rect 122104 311788 122156 311840
rect 237380 311788 237432 311840
rect 232504 309204 232556 309256
rect 237472 309204 237524 309256
rect 157248 309136 157300 309188
rect 237380 309136 237432 309188
rect 235356 307776 235408 307828
rect 237380 307776 237432 307828
rect 232596 305056 232648 305108
rect 237472 305056 237524 305108
rect 235448 304988 235500 305040
rect 237380 304988 237432 305040
rect 151728 303628 151780 303680
rect 237380 303628 237432 303680
rect 232688 302200 232740 302252
rect 237380 302200 237432 302252
rect 235540 300908 235592 300960
rect 237472 300908 237524 300960
rect 148968 300840 149020 300892
rect 237380 300840 237432 300892
rect 235632 298120 235684 298172
rect 237380 298120 237432 298172
rect 146208 296692 146260 296744
rect 237380 296692 237432 296744
rect 235724 295332 235776 295384
rect 237380 295332 237432 295384
rect 144828 293972 144880 294024
rect 237380 293972 237432 294024
rect 3148 292612 3200 292664
rect 236644 292612 236696 292664
rect 235908 292544 235960 292596
rect 237380 292544 237432 292596
rect 142068 291184 142120 291236
rect 237380 291184 237432 291236
rect 154488 290436 154540 290488
rect 238024 290436 238076 290488
rect 235172 289824 235224 289876
rect 237380 289824 237432 289876
rect 139308 288396 139360 288448
rect 237380 288396 237432 288448
rect 117228 286492 117280 286544
rect 169760 286492 169812 286544
rect 170680 286492 170732 286544
rect 192484 286492 192536 286544
rect 121368 286424 121420 286476
rect 137284 286424 137336 286476
rect 169668 286424 169720 286476
rect 192668 286424 192720 286476
rect 136548 286356 136600 286408
rect 237380 286356 237432 286408
rect 49608 286288 49660 286340
rect 180708 286288 180760 286340
rect 133788 286220 133840 286272
rect 186688 286220 186740 286272
rect 132316 286152 132368 286204
rect 186780 286152 186832 286204
rect 126888 286084 126940 286136
rect 186964 286084 187016 286136
rect 111708 286016 111760 286068
rect 191380 286016 191432 286068
rect 108948 285948 109000 286000
rect 188804 285948 188856 286000
rect 104808 285880 104860 285932
rect 187332 285880 187384 285932
rect 86868 285812 86920 285864
rect 188344 285812 188396 285864
rect 81348 285744 81400 285796
rect 196716 285744 196768 285796
rect 79968 285676 80020 285728
rect 196624 285676 196676 285728
rect 234988 285676 235040 285728
rect 237472 285676 237524 285728
rect 113824 285608 113876 285660
rect 188896 285608 188948 285660
rect 106188 285540 106240 285592
rect 188712 285540 188764 285592
rect 102048 285472 102100 285524
rect 195244 285472 195296 285524
rect 96160 285404 96212 285456
rect 193956 285404 194008 285456
rect 93676 285336 93728 285388
rect 191288 285336 191340 285388
rect 89628 285268 89680 285320
rect 189908 285268 189960 285320
rect 128728 285200 128780 285252
rect 238668 285200 238720 285252
rect 123576 285132 123628 285184
rect 238116 285132 238168 285184
rect 118608 285064 118660 285116
rect 238392 285064 238444 285116
rect 98552 284996 98604 285048
rect 238484 284996 238536 285048
rect 91192 284928 91244 284980
rect 238024 284928 238076 284980
rect 169760 284860 169812 284912
rect 238208 284860 238260 284912
rect 232872 284316 232924 284368
rect 237380 284316 237432 284368
rect 137284 283568 137336 283620
rect 238576 283568 238628 283620
rect 232780 282888 232832 282940
rect 237472 282888 237524 282940
rect 186688 282820 186740 282872
rect 237380 282820 237432 282872
rect 196808 281528 196860 281580
rect 237380 281528 237432 281580
rect 191196 280168 191248 280220
rect 237472 280168 237524 280220
rect 186780 280100 186832 280152
rect 237380 280100 237432 280152
rect 189080 278740 189132 278792
rect 192576 278740 192628 278792
rect 189816 274728 189868 274780
rect 237380 274728 237432 274780
rect 188436 274660 188488 274712
rect 237472 274660 237524 274712
rect 186964 274592 187016 274644
rect 237380 274592 237432 274644
rect 186964 271872 187016 271924
rect 237380 271872 237432 271924
rect 540336 271872 540388 271924
rect 580172 271872 580224 271924
rect 188528 269084 188580 269136
rect 237380 269084 237432 269136
rect 190000 264936 190052 264988
rect 237380 264936 237432 264988
rect 188620 262216 188672 262268
rect 237380 262216 237432 262268
rect 193864 259496 193916 259548
rect 237380 259496 237432 259548
rect 187056 259428 187108 259480
rect 237472 259428 237524 259480
rect 188896 259360 188948 259412
rect 237380 259360 237432 259412
rect 191380 256640 191432 256692
rect 237472 256640 237524 256692
rect 192760 255280 192812 255332
rect 237380 255280 237432 255332
rect 187148 253920 187200 253972
rect 237380 253920 237432 253972
rect 190092 252560 190144 252612
rect 237472 252560 237524 252612
rect 188804 252492 188856 252544
rect 237380 252492 237432 252544
rect 191380 249772 191432 249824
rect 237380 249772 237432 249824
rect 188712 248344 188764 248396
rect 237380 248344 237432 248396
rect 187240 245624 187292 245676
rect 237380 245624 237432 245676
rect 194048 244264 194100 244316
rect 237380 244264 237432 244316
rect 187332 242836 187384 242888
rect 237380 242836 237432 242888
rect 3240 240116 3292 240168
rect 46296 240116 46348 240168
rect 190184 240116 190236 240168
rect 237380 240116 237432 240168
rect 195244 237328 195296 237380
rect 237380 237328 237432 237380
rect 188712 235968 188764 236020
rect 237380 235968 237432 236020
rect 540428 231820 540480 231872
rect 580172 231820 580224 231872
rect 188804 230460 188856 230512
rect 237380 230460 237432 230512
rect 235816 227808 235868 227860
rect 237380 227808 237432 227860
rect 195244 227740 195296 227792
rect 237472 227740 237524 227792
rect 193956 227672 194008 227724
rect 237380 227672 237432 227724
rect 191472 224952 191524 225004
rect 237380 224952 237432 225004
rect 193956 223592 194008 223644
rect 237380 223592 237432 223644
rect 191288 222096 191340 222148
rect 237380 222096 237432 222148
rect 188896 220804 188948 220856
rect 237380 220804 237432 220856
rect 189080 218084 189132 218136
rect 192852 218084 192904 218136
rect 193128 218016 193180 218068
rect 237380 218016 237432 218068
rect 190276 216724 190328 216776
rect 237380 216724 237432 216776
rect 189080 216656 189132 216708
rect 191288 216656 191340 216708
rect 189172 215364 189224 215416
rect 191564 215364 191616 215416
rect 188988 215296 189040 215348
rect 237380 215296 237432 215348
rect 187332 213936 187384 213988
rect 237472 213936 237524 213988
rect 190460 213868 190512 213920
rect 237380 213868 237432 213920
rect 189080 213800 189132 213852
rect 193128 213800 193180 213852
rect 190368 212508 190420 212560
rect 237380 212508 237432 212560
rect 189908 212440 189960 212492
rect 237472 212440 237524 212492
rect 188252 209856 188304 209908
rect 237472 209856 237524 209908
rect 187424 209788 187476 209840
rect 237380 209788 237432 209840
rect 191564 209720 191616 209772
rect 237472 209720 237524 209772
rect 47584 207680 47636 207732
rect 48228 207680 48280 207732
rect 49608 207680 49660 207732
rect 189632 207000 189684 207052
rect 237380 207000 237432 207052
rect 188344 206932 188396 206984
rect 237472 206932 237524 206984
rect 188160 205640 188212 205692
rect 237380 205640 237432 205692
rect 191288 202784 191340 202836
rect 237380 202784 237432 202836
rect 189080 201492 189132 201544
rect 237380 201492 237432 201544
rect 186964 200744 187016 200796
rect 238208 200744 238260 200796
rect 188344 200132 188396 200184
rect 237380 200132 237432 200184
rect 128360 199520 128412 199572
rect 238116 199520 238168 199572
rect 120080 199452 120132 199504
rect 237840 199452 237892 199504
rect 110420 199384 110472 199436
rect 238024 199384 238076 199436
rect 111064 199316 111116 199368
rect 187148 199316 187200 199368
rect 91192 199248 91244 199300
rect 188988 199248 189040 199300
rect 88616 199180 88668 199232
rect 188252 199180 188304 199232
rect 78864 199112 78916 199164
rect 187332 199112 187384 199164
rect 77760 199044 77812 199096
rect 187424 199044 187476 199096
rect 70584 198976 70636 199028
rect 188344 198976 188396 199028
rect 103704 198908 103756 198960
rect 238576 198908 238628 198960
rect 82544 198840 82596 198892
rect 238484 198840 238536 198892
rect 80152 198772 80204 198824
rect 238300 198772 238352 198824
rect 81348 198704 81400 198756
rect 238668 198704 238720 198756
rect 86224 198636 86276 198688
rect 110420 198636 110472 198688
rect 121000 198636 121052 198688
rect 128360 198636 128412 198688
rect 105912 198568 105964 198620
rect 235632 198568 235684 198620
rect 108488 198500 108540 198552
rect 238392 198500 238444 198552
rect 71872 198432 71924 198484
rect 188160 198432 188212 198484
rect 92848 198364 92900 198416
rect 190000 198364 190052 198416
rect 93584 198296 93636 198348
rect 188896 198296 188948 198348
rect 95976 198228 96028 198280
rect 191472 198228 191524 198280
rect 98368 198160 98420 198212
rect 188804 198160 188856 198212
rect 100944 198092 100996 198144
rect 188712 198092 188764 198144
rect 106096 198024 106148 198076
rect 187240 198024 187292 198076
rect 75552 197956 75604 198008
rect 237380 197956 237432 198008
rect 113640 197888 113692 197940
rect 186964 197888 187016 197940
rect 76840 197820 76892 197872
rect 120080 197820 120132 197872
rect 123576 197820 123628 197872
rect 188528 197820 188580 197872
rect 128912 197752 128964 197804
rect 188436 197752 188488 197804
rect 47952 197684 48004 197736
rect 237932 197684 237984 197736
rect 173440 197276 173492 197328
rect 195244 197276 195296 197328
rect 48044 197208 48096 197260
rect 190276 197208 190328 197260
rect 192852 197208 192904 197260
rect 237380 197208 237432 197260
rect 85856 197140 85908 197192
rect 194048 197140 194100 197192
rect 84568 197072 84620 197124
rect 190184 197072 190236 197124
rect 87972 197004 88024 197056
rect 191380 197004 191432 197056
rect 89536 196936 89588 196988
rect 192760 196936 192812 196988
rect 90824 196868 90876 196920
rect 193864 196868 193916 196920
rect 88248 196800 88300 196852
rect 190092 196800 190144 196852
rect 118424 196732 118476 196784
rect 188620 196732 188672 196784
rect 117044 196664 117096 196716
rect 187056 196664 187108 196716
rect 73436 196596 73488 196648
rect 238024 196596 238076 196648
rect 126612 196528 126664 196580
rect 186872 196528 186924 196580
rect 83648 196460 83700 196512
rect 237472 196460 237524 196512
rect 173256 196392 173308 196444
rect 193956 196392 194008 196444
rect 49516 195916 49568 195968
rect 237380 195916 237432 195968
rect 69664 195848 69716 195900
rect 237472 195848 237524 195900
rect 107016 195780 107068 195832
rect 235540 195780 235592 195832
rect 108580 195712 108632 195764
rect 235448 195712 235500 195764
rect 109224 195644 109276 195696
rect 235356 195644 235408 195696
rect 138664 195576 138716 195628
rect 237104 195576 237156 195628
rect 141240 195508 141292 195560
rect 237012 195508 237064 195560
rect 143448 195440 143500 195492
rect 236920 195440 236972 195492
rect 146024 195372 146076 195424
rect 236828 195372 236880 195424
rect 148600 195304 148652 195356
rect 236736 195304 236788 195356
rect 150992 195236 151044 195288
rect 232688 195236 232740 195288
rect 153384 195168 153436 195220
rect 232596 195168 232648 195220
rect 133512 195100 133564 195152
rect 196808 195100 196860 195152
rect 155960 194488 156012 194540
rect 232504 194488 232556 194540
rect 196716 194420 196768 194472
rect 237380 194420 237432 194472
rect 81256 193128 81308 193180
rect 237380 193128 237432 193180
rect 74356 191768 74408 191820
rect 237380 191768 237432 191820
rect 192668 191700 192720 191752
rect 237472 191700 237524 191752
rect 67548 190408 67600 190460
rect 237380 190408 237432 190460
rect 68928 188980 68980 189032
rect 238392 188980 238444 189032
rect 3332 187688 3384 187740
rect 239128 187688 239180 187740
rect 78588 187620 78640 187672
rect 238760 187620 238812 187672
rect 196624 187552 196676 187604
rect 238392 187552 238444 187604
rect 192484 184832 192536 184884
rect 238760 184832 238812 184884
rect 49332 183472 49384 183524
rect 238300 183472 238352 183524
rect 66168 183404 66220 183456
rect 238392 183404 238444 183456
rect 239036 182860 239088 182912
rect 239680 182860 239732 182912
rect 239312 182724 239364 182776
rect 239680 182724 239732 182776
rect 192576 182112 192628 182164
rect 239404 182112 239456 182164
rect 49424 181432 49476 181484
rect 238576 181432 238628 181484
rect 47584 181296 47636 181348
rect 48228 181296 48280 181348
rect 48228 180820 48280 180872
rect 87972 180820 88024 180872
rect 300216 180208 300268 180260
rect 580172 180208 580224 180260
rect 300124 180140 300176 180192
rect 580908 180140 580960 180192
rect 297916 179868 297968 179920
rect 580816 180072 580868 180124
rect 390192 179664 390244 179716
rect 538312 179664 538364 179716
rect 318248 179596 318300 179648
rect 540244 179596 540296 179648
rect 310336 179528 310388 179580
rect 540336 179528 540388 179580
rect 302240 179460 302292 179512
rect 540428 179460 540480 179512
rect 338028 179392 338080 179444
rect 577504 179392 577556 179444
rect 46296 179324 46348 179376
rect 517612 179324 517664 179376
rect 44824 179256 44876 179308
rect 493600 179256 493652 179308
rect 46204 179188 46256 179240
rect 485780 179188 485832 179240
rect 239128 179120 239180 179172
rect 521660 179120 521712 179172
rect 236644 179052 236696 179104
rect 509608 179052 509660 179104
rect 536932 179052 536984 179104
rect 538404 179052 538456 179104
rect 233884 178984 233936 179036
rect 501604 178984 501656 179036
rect 191104 178916 191156 178968
rect 449992 178916 450044 178968
rect 239496 178848 239548 178900
rect 477592 178848 477644 178900
rect 239864 178780 239916 178832
rect 280068 178780 280120 178832
rect 355692 178780 355744 178832
rect 580724 178780 580776 178832
rect 239220 178712 239272 178764
rect 282920 178712 282972 178764
rect 310428 178712 310480 178764
rect 580080 178712 580132 178764
rect 3700 178644 3752 178696
rect 401600 178644 401652 178696
rect 408500 178644 408552 178696
rect 580632 178644 580684 178696
rect 189724 178576 189776 178628
rect 410064 178576 410116 178628
rect 366272 178508 366324 178560
rect 580264 178508 580316 178560
rect 239680 178440 239732 178492
rect 393596 178440 393648 178492
rect 406200 178032 406252 178084
rect 580172 178032 580224 178084
rect 334256 177964 334308 178016
rect 355692 177964 355744 178016
rect 531964 177964 532016 178016
rect 538036 177964 538088 178016
rect 289912 177896 289964 177948
rect 300124 177896 300176 177948
rect 3884 177828 3936 177880
rect 490012 177828 490064 177880
rect 3792 177760 3844 177812
rect 481640 177760 481692 177812
rect 490564 177760 490616 177812
rect 513564 177760 513616 177812
rect 530676 177760 530728 177812
rect 536932 177760 536984 177812
rect 87972 177692 88024 177744
rect 241980 177692 242032 177744
rect 281908 177692 281960 177744
rect 300216 177692 300268 177744
rect 342168 177692 342220 177744
rect 580540 177692 580592 177744
rect 306196 177624 306248 177676
rect 538956 177624 539008 177676
rect 293960 177556 294012 177608
rect 310428 177556 310480 177608
rect 350264 177556 350316 177608
rect 580448 177556 580500 177608
rect 314200 177488 314252 177540
rect 538864 177488 538916 177540
rect 358176 177420 358228 177472
rect 580356 177420 580408 177472
rect 362224 177352 362276 177404
rect 542360 177352 542412 177404
rect 1400 177284 1452 177336
rect 245936 177284 245988 177336
rect 382188 177284 382240 177336
rect 538220 177284 538272 177336
rect 239036 177216 239088 177268
rect 413560 177216 413612 177268
rect 273904 177148 273956 177200
rect 406200 177148 406252 177200
rect 322296 177080 322348 177132
rect 408500 177080 408552 177132
rect 4068 177012 4120 177064
rect 505560 177012 505612 177064
rect 3976 176944 4028 176996
rect 497556 176944 497608 176996
rect 3516 176604 3568 176656
rect 461584 176604 461636 176656
rect 23480 176536 23532 176588
rect 425612 176536 425664 176588
rect 330208 176468 330260 176520
rect 577596 176468 577648 176520
rect 326344 176400 326396 176452
rect 543004 176400 543056 176452
rect 378048 176332 378100 176384
rect 531964 176332 532016 176384
rect 282920 176264 282972 176316
rect 385592 176264 385644 176316
rect 398288 176264 398340 176316
rect 530676 176264 530728 176316
rect 280068 176196 280120 176248
rect 405740 176196 405792 176248
rect 235264 175176 235316 175228
rect 457536 175176 457588 175228
rect 256700 174088 256752 174140
rect 257896 174088 257948 174140
rect 285680 153144 285732 153196
rect 580172 153144 580224 153196
rect 3424 150356 3476 150408
rect 490564 150356 490616 150408
rect 264980 139340 265032 139392
rect 580172 139340 580224 139392
rect 3240 137912 3292 137964
rect 525800 137912 525852 137964
rect 277400 113092 277452 113144
rect 579804 113092 579856 113144
rect 256700 100648 256752 100700
rect 580172 100648 580224 100700
rect 3148 85484 3200 85536
rect 529940 85484 529992 85536
rect 269120 73108 269172 73160
rect 580172 73108 580224 73160
rect 249800 60664 249852 60716
rect 580172 60664 580224 60716
rect 3424 45500 3476 45552
rect 532700 45500 532752 45552
rect 260840 33056 260892 33108
rect 580172 33056 580224 33108
rect 3424 6808 3476 6860
rect 536840 6808 536892 6860
rect 253940 6740 253992 6792
rect 580172 6740 580224 6792
rect 572 3408 624 3460
rect 47584 3408 47636 3460
<< metal2 >>
rect 8086 703520 8198 704960
rect 23492 703582 24164 703610
rect 8128 700369 8156 703520
rect 8114 700360 8170 700369
rect 8114 700295 8170 700304
rect 3422 671256 3478 671265
rect 3422 671191 3478 671200
rect 3054 566944 3110 566953
rect 3054 566879 3110 566888
rect 3068 565894 3096 566879
rect 3056 565888 3108 565894
rect 3056 565830 3108 565836
rect 3330 514856 3386 514865
rect 3330 514791 3332 514800
rect 3384 514791 3386 514800
rect 3332 514762 3384 514768
rect 3330 501800 3386 501809
rect 3330 501735 3386 501744
rect 3344 501022 3372 501735
rect 3332 501016 3384 501022
rect 3332 500958 3384 500964
rect 3330 449576 3386 449585
rect 3330 449511 3386 449520
rect 3344 448594 3372 449511
rect 3332 448588 3384 448594
rect 3332 448530 3384 448536
rect 3332 397520 3384 397526
rect 3330 397488 3332 397497
rect 3384 397488 3386 397497
rect 3330 397423 3386 397432
rect 3054 345400 3110 345409
rect 3054 345335 3110 345344
rect 3068 345098 3096 345335
rect 3056 345092 3108 345098
rect 3056 345034 3108 345040
rect 3146 293176 3202 293185
rect 3146 293111 3202 293120
rect 3160 292670 3188 293111
rect 3148 292664 3200 292670
rect 3148 292606 3200 292612
rect 3238 241088 3294 241097
rect 3238 241023 3294 241032
rect 3252 240174 3280 241023
rect 3240 240168 3292 240174
rect 3240 240110 3292 240116
rect 3330 188864 3386 188873
rect 3330 188799 3386 188808
rect 3344 187746 3372 188799
rect 3332 187740 3384 187746
rect 3332 187682 3384 187688
rect 3436 177857 3464 671191
rect 3514 658200 3570 658209
rect 3514 658135 3570 658144
rect 3528 656946 3556 658135
rect 3516 656940 3568 656946
rect 3516 656882 3568 656888
rect 3514 606112 3570 606121
rect 3514 606047 3570 606056
rect 3422 177848 3478 177857
rect 3422 177783 3478 177792
rect 1400 177336 1452 177342
rect 1400 177278 1452 177284
rect 572 3460 624 3466
rect 572 3402 624 3408
rect 584 480 612 3402
rect 542 -960 654 480
rect 1412 354 1440 177278
rect 3528 176662 3556 606047
rect 3606 553888 3662 553897
rect 3606 553823 3662 553832
rect 3620 553450 3648 553823
rect 3608 553444 3660 553450
rect 3608 553386 3660 553392
rect 3606 462632 3662 462641
rect 3606 462567 3662 462576
rect 3620 177993 3648 462567
rect 3698 410544 3754 410553
rect 3698 410479 3754 410488
rect 3712 178702 3740 410479
rect 3790 358456 3846 358465
rect 3790 358391 3846 358400
rect 3700 178696 3752 178702
rect 3700 178638 3752 178644
rect 3606 177984 3662 177993
rect 3606 177919 3662 177928
rect 3804 177818 3832 358391
rect 3882 306232 3938 306241
rect 3882 306167 3938 306176
rect 3896 177886 3924 306167
rect 3974 254144 4030 254153
rect 3974 254079 4030 254088
rect 3884 177880 3936 177886
rect 3884 177822 3936 177828
rect 3792 177812 3844 177818
rect 3792 177754 3844 177760
rect 3988 177002 4016 254079
rect 4066 201920 4122 201929
rect 4066 201855 4122 201864
rect 4080 177070 4108 201855
rect 4068 177064 4120 177070
rect 4068 177006 4120 177012
rect 3976 176996 4028 177002
rect 3976 176938 4028 176944
rect 3516 176656 3568 176662
rect 3516 176598 3568 176604
rect 23492 176594 23520 703582
rect 24136 703474 24164 703582
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218072 703582 218836 703610
rect 24320 703474 24348 703520
rect 24136 703446 24348 703474
rect 72988 700330 73016 703520
rect 89180 700505 89208 703520
rect 137848 700641 137876 703520
rect 137834 700632 137890 700641
rect 137834 700567 137890 700576
rect 89166 700496 89222 700505
rect 89166 700431 89222 700440
rect 154132 700398 154160 703520
rect 202800 703050 202828 703520
rect 201500 703044 201552 703050
rect 201500 702986 201552 702992
rect 202788 703044 202840 703050
rect 202788 702986 202840 702992
rect 154120 700392 154172 700398
rect 154120 700334 154172 700340
rect 189724 700392 189776 700398
rect 189724 700334 189776 700340
rect 72976 700324 73028 700330
rect 72976 700266 73028 700272
rect 157248 478916 157300 478922
rect 157248 478858 157300 478864
rect 154488 473408 154540 473414
rect 154488 473350 154540 473356
rect 151360 469260 151412 469266
rect 151360 469202 151412 469208
rect 151372 466313 151400 469202
rect 151358 466304 151414 466313
rect 151358 466239 151414 466248
rect 146024 465860 146076 465866
rect 146024 465802 146076 465808
rect 141056 465792 141108 465798
rect 141056 465734 141108 465740
rect 136088 465724 136140 465730
rect 136088 465666 136140 465672
rect 128728 465656 128780 465662
rect 128728 465598 128780 465604
rect 111064 465588 111116 465594
rect 111064 465530 111116 465536
rect 108488 465520 108540 465526
rect 108488 465462 108540 465468
rect 101312 465452 101364 465458
rect 101312 465394 101364 465400
rect 96160 465248 96212 465254
rect 91190 465216 91246 465225
rect 91190 465151 91246 465160
rect 93674 465216 93730 465225
rect 93674 465151 93676 465160
rect 91204 465118 91232 465151
rect 93728 465151 93730 465160
rect 96158 465216 96160 465225
rect 101324 465225 101352 465394
rect 106188 465384 106240 465390
rect 106188 465326 106240 465332
rect 103704 465316 103756 465322
rect 103704 465258 103756 465264
rect 103716 465225 103744 465258
rect 106200 465225 106228 465326
rect 108500 465225 108528 465462
rect 111076 465225 111104 465530
rect 128740 465225 128768 465598
rect 136100 465225 136128 465666
rect 141068 465225 141096 465734
rect 146036 465225 146064 465802
rect 154500 465225 154528 473350
rect 157260 466449 157288 478858
rect 157246 466440 157302 466449
rect 157246 466375 157302 466384
rect 169760 465996 169812 466002
rect 169760 465938 169812 465944
rect 168472 465928 168524 465934
rect 168472 465870 168524 465876
rect 168484 465225 168512 465870
rect 169772 465225 169800 465938
rect 186688 465860 186740 465866
rect 186688 465802 186740 465808
rect 96212 465216 96214 465225
rect 96158 465151 96214 465160
rect 101310 465216 101366 465225
rect 101310 465151 101366 465160
rect 103702 465216 103758 465225
rect 103702 465151 103758 465160
rect 106186 465216 106242 465225
rect 106186 465151 106242 465160
rect 108486 465216 108542 465225
rect 108486 465151 108542 465160
rect 111062 465216 111118 465225
rect 111062 465151 111118 465160
rect 128726 465216 128782 465225
rect 128726 465151 128782 465160
rect 136086 465216 136142 465225
rect 136086 465151 136142 465160
rect 141054 465216 141110 465225
rect 141054 465151 141110 465160
rect 146022 465216 146078 465225
rect 146022 465151 146078 465160
rect 154486 465216 154542 465225
rect 154486 465151 154542 465160
rect 168470 465216 168526 465225
rect 168470 465151 168526 465160
rect 169758 465216 169814 465225
rect 169758 465151 169814 465160
rect 93676 465122 93728 465128
rect 91192 465112 91244 465118
rect 91192 465054 91244 465060
rect 148508 465044 148560 465050
rect 148508 464986 148560 464992
rect 121000 464976 121052 464982
rect 121000 464918 121052 464924
rect 98552 464840 98604 464846
rect 98552 464782 98604 464788
rect 88524 464636 88576 464642
rect 88524 464578 88576 464584
rect 83464 464568 83516 464574
rect 83464 464510 83516 464516
rect 83476 463729 83504 464510
rect 88536 463729 88564 464578
rect 98564 463729 98592 464782
rect 118608 464500 118660 464506
rect 118608 464442 118660 464448
rect 116124 464432 116176 464438
rect 116124 464374 116176 464380
rect 113640 464364 113692 464370
rect 113640 464306 113692 464312
rect 113652 463729 113680 464306
rect 116136 463729 116164 464374
rect 118620 463729 118648 464442
rect 121012 463729 121040 464918
rect 143632 464908 143684 464914
rect 143632 464850 143684 464856
rect 133512 464772 133564 464778
rect 133512 464714 133564 464720
rect 131120 464704 131172 464710
rect 131120 464646 131172 464652
rect 123576 464296 123628 464302
rect 123576 464238 123628 464244
rect 123588 463729 123616 464238
rect 125968 464228 126020 464234
rect 125968 464170 126020 464176
rect 125980 463729 126008 464170
rect 131132 464001 131160 464646
rect 131118 463992 131174 464001
rect 131118 463927 131174 463936
rect 133524 463729 133552 464714
rect 138480 464160 138532 464166
rect 138480 464102 138532 464108
rect 138492 463729 138520 464102
rect 143644 463729 143672 464850
rect 148520 463729 148548 464986
rect 83462 463720 83518 463729
rect 83462 463655 83518 463664
rect 88522 463720 88578 463729
rect 88522 463655 88578 463664
rect 98550 463720 98606 463729
rect 98550 463655 98606 463664
rect 113638 463720 113694 463729
rect 113638 463655 113694 463664
rect 116122 463720 116178 463729
rect 116122 463655 116178 463664
rect 118606 463720 118662 463729
rect 118606 463655 118662 463664
rect 120998 463720 121054 463729
rect 120998 463655 121054 463664
rect 123574 463720 123630 463729
rect 123574 463655 123630 463664
rect 125966 463720 126022 463729
rect 125966 463655 126022 463664
rect 133510 463720 133566 463729
rect 133510 463655 133566 463664
rect 138478 463720 138534 463729
rect 138478 463655 138534 463664
rect 143630 463720 143686 463729
rect 143630 463655 143686 463664
rect 148506 463720 148562 463729
rect 148506 463655 148562 463664
rect 186700 463010 186728 465802
rect 187240 465792 187292 465798
rect 187240 465734 187292 465740
rect 187148 465724 187200 465730
rect 187148 465666 187200 465672
rect 187056 465656 187108 465662
rect 187056 465598 187108 465604
rect 186964 465588 187016 465594
rect 186964 465530 187016 465536
rect 186688 463004 186740 463010
rect 186688 462946 186740 462952
rect 46204 448588 46256 448594
rect 46204 448530 46256 448536
rect 44824 397520 44876 397526
rect 44824 397462 44876 397468
rect 44836 179314 44864 397462
rect 44824 179308 44876 179314
rect 44824 179250 44876 179256
rect 46216 179246 46244 448530
rect 48042 416936 48098 416945
rect 48042 416871 48098 416880
rect 47950 415984 48006 415993
rect 47950 415919 48006 415928
rect 47582 388376 47638 388385
rect 47582 388311 47638 388320
rect 46296 240168 46348 240174
rect 46296 240110 46348 240116
rect 46308 179382 46336 240110
rect 47596 207738 47624 388311
rect 47858 388104 47914 388113
rect 47858 388039 47914 388048
rect 47872 371890 47900 388039
rect 47860 371884 47912 371890
rect 47860 371826 47912 371832
rect 47964 369170 47992 415919
rect 47952 369164 48004 369170
rect 47952 369106 48004 369112
rect 48056 358766 48084 416871
rect 48226 413808 48282 413817
rect 48226 413743 48282 413752
rect 48134 390008 48190 390017
rect 48134 389943 48190 389952
rect 48044 358760 48096 358766
rect 48044 358702 48096 358708
rect 48148 313274 48176 389943
rect 48240 379574 48268 413743
rect 49330 412856 49386 412865
rect 49330 412791 49386 412800
rect 49238 410000 49294 410009
rect 49238 409935 49294 409944
rect 48228 379568 48280 379574
rect 48228 379510 48280 379516
rect 49252 332586 49280 409935
rect 49344 376038 49372 412791
rect 49422 411074 49478 411083
rect 49422 411009 49478 411018
rect 49332 376032 49384 376038
rect 49332 375974 49384 375980
rect 49436 365022 49464 411009
rect 49606 408218 49662 408227
rect 49606 408153 49662 408162
rect 49424 365016 49476 365022
rect 49424 364958 49476 364964
rect 49240 332580 49292 332586
rect 49240 332522 49292 332528
rect 49620 327078 49648 408153
rect 186976 389162 187004 465530
rect 187068 423638 187096 465598
rect 187160 440230 187188 465666
rect 187252 449886 187280 465734
rect 188344 465520 188396 465526
rect 188344 465462 188396 465468
rect 187240 449880 187292 449886
rect 187240 449822 187292 449828
rect 187148 440224 187200 440230
rect 187148 440166 187200 440172
rect 187056 423632 187108 423638
rect 187056 423574 187108 423580
rect 187056 416832 187108 416838
rect 187056 416774 187108 416780
rect 186964 389156 187016 389162
rect 186964 389098 187016 389104
rect 186964 386436 187016 386442
rect 186964 386378 187016 386384
rect 186688 380180 186740 380186
rect 186688 380122 186740 380128
rect 110970 379672 111026 379681
rect 110970 379607 111026 379616
rect 113546 379672 113602 379681
rect 113546 379607 113602 379616
rect 118330 379672 118386 379681
rect 118330 379607 118386 379616
rect 120998 379672 121054 379681
rect 120998 379607 121054 379616
rect 123482 379672 123538 379681
rect 123482 379607 123538 379616
rect 130934 379672 130990 379681
rect 130934 379607 130990 379616
rect 144918 379672 144974 379681
rect 144918 379607 144974 379616
rect 49884 379568 49936 379574
rect 49884 379510 49936 379516
rect 87050 379536 87106 379545
rect 49896 349110 49924 379510
rect 87050 379471 87106 379480
rect 88154 379536 88210 379545
rect 88154 379471 88210 379480
rect 89442 379536 89498 379545
rect 89442 379471 89498 379480
rect 90730 379536 90786 379545
rect 90730 379471 90786 379480
rect 87064 378962 87092 379471
rect 88168 379098 88196 379471
rect 89456 379166 89484 379471
rect 89444 379160 89496 379166
rect 89444 379102 89496 379108
rect 88156 379092 88208 379098
rect 88156 379034 88208 379040
rect 90744 379030 90772 379471
rect 110984 379370 111012 379607
rect 113560 379438 113588 379607
rect 116030 379536 116086 379545
rect 116030 379471 116032 379480
rect 116084 379471 116086 379480
rect 116032 379442 116084 379448
rect 113548 379432 113600 379438
rect 113548 379374 113600 379380
rect 110972 379364 111024 379370
rect 110972 379306 111024 379312
rect 90732 379024 90784 379030
rect 90732 378966 90784 378972
rect 87052 378956 87104 378962
rect 87052 378898 87104 378904
rect 118344 378758 118372 379607
rect 121012 378826 121040 379607
rect 121000 378820 121052 378826
rect 121000 378762 121052 378768
rect 118332 378752 118384 378758
rect 118332 378694 118384 378700
rect 123496 378690 123524 379607
rect 123484 378684 123536 378690
rect 123484 378626 123536 378632
rect 130948 378622 130976 379607
rect 144932 379234 144960 379607
rect 150990 379536 151046 379545
rect 150990 379471 151046 379480
rect 151004 379302 151032 379471
rect 150992 379296 151044 379302
rect 150992 379238 151044 379244
rect 144920 379228 144972 379234
rect 144920 379170 144972 379176
rect 135996 378888 136048 378894
rect 135996 378830 136048 378836
rect 130936 378616 130988 378622
rect 130936 378558 130988 378564
rect 91928 378072 91980 378078
rect 67546 378040 67602 378049
rect 67546 377975 67602 377984
rect 74354 378040 74410 378049
rect 74354 377975 74410 377984
rect 78494 378040 78550 378049
rect 78494 377975 78550 377984
rect 81162 378040 81218 378049
rect 81162 377975 81218 377984
rect 85946 378040 86002 378049
rect 85946 377975 86002 377984
rect 91926 378040 91928 378049
rect 91980 378040 91982 378049
rect 91926 377975 91982 377984
rect 92846 378040 92902 378049
rect 92846 377975 92848 377984
rect 66166 377088 66222 377097
rect 66166 377023 66222 377032
rect 49884 349104 49936 349110
rect 49884 349046 49936 349052
rect 49608 327072 49660 327078
rect 49608 327014 49660 327020
rect 66180 314634 66208 377023
rect 67560 321570 67588 377975
rect 68926 377088 68982 377097
rect 68926 377023 68982 377032
rect 70306 377088 70362 377097
rect 70306 377023 70362 377032
rect 71686 377088 71742 377097
rect 71686 377023 71742 377032
rect 73066 377088 73122 377097
rect 73066 377023 73122 377032
rect 67548 321564 67600 321570
rect 67548 321506 67600 321512
rect 68940 320142 68968 377023
rect 70320 325650 70348 377023
rect 71700 332518 71728 377023
rect 73080 338094 73108 377023
rect 73068 338088 73120 338094
rect 73068 338030 73120 338036
rect 71688 332512 71740 332518
rect 71688 332454 71740 332460
rect 70308 325644 70360 325650
rect 70308 325586 70360 325592
rect 74368 324970 74396 377975
rect 75826 377088 75882 377097
rect 75826 377023 75882 377032
rect 77206 377088 77262 377097
rect 77206 377023 77262 377032
rect 78310 377088 78366 377097
rect 78310 377023 78312 377032
rect 74446 376952 74502 376961
rect 74446 376887 74502 376896
rect 74356 324964 74408 324970
rect 74356 324906 74408 324912
rect 74460 323610 74488 376887
rect 75840 329798 75868 377023
rect 77220 335306 77248 377023
rect 78364 377023 78366 377032
rect 78312 376994 78364 377000
rect 78508 340882 78536 377975
rect 79966 377088 80022 377097
rect 79324 377052 79376 377058
rect 79966 377023 80022 377032
rect 79324 376994 79376 377000
rect 78496 340876 78548 340882
rect 78496 340818 78548 340824
rect 77208 335300 77260 335306
rect 77208 335242 77260 335248
rect 75828 329792 75880 329798
rect 75828 329734 75880 329740
rect 74448 323604 74500 323610
rect 74448 323546 74500 323552
rect 68928 320136 68980 320142
rect 68928 320078 68980 320084
rect 79336 317422 79364 376994
rect 79980 346390 80008 377023
rect 81176 356046 81204 377975
rect 81254 377088 81310 377097
rect 81254 377023 81310 377032
rect 82726 377088 82782 377097
rect 82726 377023 82782 377032
rect 84106 377088 84162 377097
rect 84106 377023 84162 377032
rect 85486 377088 85542 377097
rect 85486 377023 85542 377032
rect 81164 356040 81216 356046
rect 81164 355982 81216 355988
rect 81268 351898 81296 377023
rect 81346 376952 81402 376961
rect 81346 376887 81402 376896
rect 81256 351892 81308 351898
rect 81256 351834 81308 351840
rect 79968 346384 80020 346390
rect 79968 346326 80020 346332
rect 81360 324290 81388 376887
rect 82740 361554 82768 377023
rect 84014 376952 84070 376961
rect 84014 376887 84070 376896
rect 84028 367062 84056 376887
rect 84016 367056 84068 367062
rect 84016 366998 84068 367004
rect 82728 361548 82780 361554
rect 82728 361490 82780 361496
rect 84120 329730 84148 377023
rect 85500 371210 85528 377023
rect 85960 376718 85988 377975
rect 92900 377975 92902 377984
rect 93950 378040 94006 378049
rect 93950 377975 94006 377984
rect 95238 378040 95294 378049
rect 95238 377975 95294 377984
rect 96526 378040 96582 378049
rect 96526 377975 96582 377984
rect 97630 378040 97686 378049
rect 97630 377975 97686 377984
rect 99930 378040 99986 378049
rect 99930 377975 99986 377984
rect 104806 378040 104862 378049
rect 104806 377975 104862 377984
rect 106094 378040 106150 378049
rect 106094 377975 106150 377984
rect 108486 378040 108542 378049
rect 108486 377975 108542 377984
rect 125966 378040 126022 378049
rect 125966 377975 126022 377984
rect 128542 378040 128598 378049
rect 128542 377975 128598 377984
rect 133510 378040 133566 378049
rect 133510 377975 133566 377984
rect 92848 377946 92900 377952
rect 93964 377942 93992 377975
rect 93952 377936 94004 377942
rect 93952 377878 94004 377884
rect 95252 377874 95280 377975
rect 96434 377904 96490 377913
rect 95240 377868 95292 377874
rect 96434 377839 96490 377848
rect 95240 377810 95292 377816
rect 96448 377806 96476 377839
rect 96436 377800 96488 377806
rect 96436 377742 96488 377748
rect 86774 377088 86830 377097
rect 86774 377023 86830 377032
rect 89626 377088 89682 377097
rect 89626 377023 89682 377032
rect 92386 377088 92442 377097
rect 92386 377023 92442 377032
rect 93766 377088 93822 377097
rect 93766 377023 93822 377032
rect 85948 376712 86000 376718
rect 85948 376654 86000 376660
rect 85488 371204 85540 371210
rect 85488 371146 85540 371152
rect 86788 336734 86816 377023
rect 89640 342242 89668 377023
rect 92400 347750 92428 377023
rect 93780 351830 93808 377023
rect 96540 357406 96568 377975
rect 97644 376650 97672 377975
rect 99944 377194 99972 377975
rect 102046 377768 102102 377777
rect 102046 377703 102102 377712
rect 99932 377188 99984 377194
rect 99932 377130 99984 377136
rect 99286 377088 99342 377097
rect 99286 377023 99342 377032
rect 97632 376644 97684 376650
rect 97632 376586 97684 376592
rect 99300 362914 99328 377023
rect 102060 366994 102088 377703
rect 104820 372570 104848 377975
rect 106108 377466 106136 377975
rect 108500 377534 108528 377975
rect 125980 377738 126008 377975
rect 125968 377732 126020 377738
rect 125968 377674 126020 377680
rect 128556 377670 128584 377975
rect 128544 377664 128596 377670
rect 128544 377606 128596 377612
rect 133524 377602 133552 377975
rect 133512 377596 133564 377602
rect 133512 377538 133564 377544
rect 136008 377534 136036 378830
rect 140778 378720 140834 378729
rect 140778 378655 140834 378664
rect 136086 378040 136142 378049
rect 136086 377975 136142 377984
rect 138662 378040 138718 378049
rect 138662 377975 138718 377984
rect 136100 377534 136128 377975
rect 108488 377528 108540 377534
rect 108488 377470 108540 377476
rect 135996 377528 136048 377534
rect 135996 377470 136048 377476
rect 136088 377528 136140 377534
rect 136088 377470 136140 377476
rect 106096 377460 106148 377466
rect 106096 377402 106148 377408
rect 138676 377398 138704 377975
rect 140792 377806 140820 378655
rect 141146 378040 141202 378049
rect 141146 377975 141202 377984
rect 146022 378040 146078 378049
rect 146022 377975 146078 377984
rect 148598 378040 148654 378049
rect 148598 377975 148654 377984
rect 153382 378040 153438 378049
rect 153382 377975 153438 377984
rect 155958 378040 156014 378049
rect 155958 377975 156014 377984
rect 140780 377800 140832 377806
rect 140780 377742 140832 377748
rect 138664 377392 138716 377398
rect 138664 377334 138716 377340
rect 141160 377330 141188 377975
rect 141148 377324 141200 377330
rect 141148 377266 141200 377272
rect 146036 377262 146064 377975
rect 148612 377806 148640 377975
rect 148600 377800 148652 377806
rect 148600 377742 148652 377748
rect 146024 377256 146076 377262
rect 146024 377198 146076 377204
rect 153396 376582 153424 377975
rect 153384 376576 153436 376582
rect 153384 376518 153436 376524
rect 155972 376514 156000 377975
rect 186700 377942 186728 380122
rect 186976 379370 187004 386378
rect 186964 379364 187016 379370
rect 186964 379306 187016 379312
rect 186688 377936 186740 377942
rect 186688 377878 186740 377884
rect 187068 377738 187096 416774
rect 187148 415472 187200 415478
rect 187148 415414 187200 415420
rect 187160 377874 187188 415414
rect 187240 411324 187292 411330
rect 187240 411266 187292 411272
rect 187252 378690 187280 411266
rect 187332 401668 187384 401674
rect 187332 401610 187384 401616
rect 187344 378758 187372 401610
rect 187424 396092 187476 396098
rect 187424 396034 187476 396040
rect 187436 379506 187464 396034
rect 187516 392012 187568 392018
rect 187516 391954 187568 391960
rect 187424 379500 187476 379506
rect 187424 379442 187476 379448
rect 187528 379438 187556 391954
rect 188252 390584 188304 390590
rect 188252 390526 188304 390532
rect 187792 385076 187844 385082
rect 187792 385018 187844 385024
rect 187700 380928 187752 380934
rect 187700 380870 187752 380876
rect 187516 379432 187568 379438
rect 187516 379374 187568 379380
rect 187712 378962 187740 380870
rect 187804 379098 187832 385018
rect 188264 379166 188292 390526
rect 188356 383654 188384 465462
rect 188620 464160 188672 464166
rect 188620 464102 188672 464108
rect 188436 458244 188488 458250
rect 188436 458186 188488 458192
rect 188344 383648 188396 383654
rect 188344 383590 188396 383596
rect 188252 379160 188304 379166
rect 188252 379102 188304 379108
rect 187792 379092 187844 379098
rect 187792 379034 187844 379040
rect 187700 378956 187752 378962
rect 187700 378898 187752 378904
rect 187332 378752 187384 378758
rect 187332 378694 187384 378700
rect 187240 378684 187292 378690
rect 187240 378626 187292 378632
rect 187148 377868 187200 377874
rect 187148 377810 187200 377816
rect 187056 377732 187108 377738
rect 187056 377674 187108 377680
rect 180706 377360 180762 377369
rect 180706 377295 180762 377304
rect 173806 377224 173862 377233
rect 173806 377159 173862 377168
rect 173714 376952 173770 376961
rect 173714 376887 173770 376896
rect 155960 376508 156012 376514
rect 155960 376450 156012 376456
rect 104808 372564 104860 372570
rect 104808 372506 104860 372512
rect 122104 371884 122156 371890
rect 122104 371826 122156 371832
rect 102048 366988 102100 366994
rect 102048 366930 102100 366936
rect 99288 362908 99340 362914
rect 99288 362850 99340 362856
rect 96528 357400 96580 357406
rect 96528 357342 96580 357348
rect 93768 351824 93820 351830
rect 93768 351766 93820 351772
rect 92388 347744 92440 347750
rect 92388 347686 92440 347692
rect 89628 342236 89680 342242
rect 89628 342178 89680 342184
rect 86776 336728 86828 336734
rect 86776 336670 86828 336676
rect 84108 329724 84160 329730
rect 84108 329666 84160 329672
rect 81348 324284 81400 324290
rect 81348 324226 81400 324232
rect 79324 317416 79376 317422
rect 79324 317358 79376 317364
rect 66168 314628 66220 314634
rect 66168 314570 66220 314576
rect 48136 313268 48188 313274
rect 48136 313210 48188 313216
rect 122116 311846 122144 371826
rect 173728 360194 173756 376887
rect 173716 360188 173768 360194
rect 173716 360130 173768 360136
rect 173820 355978 173848 377159
rect 177304 369164 177356 369170
rect 177304 369106 177356 369112
rect 173808 355972 173860 355978
rect 173808 355914 173860 355920
rect 177316 354686 177344 369106
rect 177304 354680 177356 354686
rect 177304 354622 177356 354628
rect 122104 311840 122156 311846
rect 122104 311782 122156 311788
rect 157248 309188 157300 309194
rect 157248 309130 157300 309136
rect 151728 303680 151780 303686
rect 151728 303622 151780 303628
rect 148968 300892 149020 300898
rect 148968 300834 149020 300840
rect 146208 296744 146260 296750
rect 146208 296686 146260 296692
rect 144828 294024 144880 294030
rect 144828 293966 144880 293972
rect 142068 291236 142120 291242
rect 142068 291178 142120 291184
rect 139308 288448 139360 288454
rect 139308 288390 139360 288396
rect 117228 286544 117280 286550
rect 117226 286512 117228 286521
rect 117280 286512 117282 286521
rect 117226 286447 117282 286456
rect 121368 286476 121420 286482
rect 121368 286418 121420 286424
rect 137284 286476 137336 286482
rect 137284 286418 137336 286424
rect 49608 286340 49660 286346
rect 49608 286282 49660 286288
rect 48134 236872 48190 236881
rect 48134 236807 48190 236816
rect 47950 235920 48006 235929
rect 47950 235855 48006 235864
rect 47766 232792 47822 232801
rect 47766 232727 47822 232736
rect 47674 231024 47730 231033
rect 47674 230959 47730 230968
rect 47584 207732 47636 207738
rect 47584 207674 47636 207680
rect 47688 199617 47716 230959
rect 47780 199753 47808 232727
rect 47858 229936 47914 229945
rect 47858 229871 47914 229880
rect 47766 199744 47822 199753
rect 47766 199679 47822 199688
rect 47674 199608 47730 199617
rect 47674 199543 47730 199552
rect 47872 197305 47900 229871
rect 47964 197742 47992 235855
rect 48042 233744 48098 233753
rect 48042 233679 48098 233688
rect 47952 197736 48004 197742
rect 47952 197678 48004 197684
rect 47858 197296 47914 197305
rect 48056 197266 48084 233679
rect 48148 199889 48176 236807
rect 49514 228218 49570 228227
rect 49514 228153 49570 228162
rect 49330 209944 49386 209953
rect 49330 209879 49386 209888
rect 48228 207732 48280 207738
rect 48228 207674 48280 207680
rect 48134 199880 48190 199889
rect 48134 199815 48190 199824
rect 47858 197231 47914 197240
rect 48044 197260 48096 197266
rect 48044 197202 48096 197208
rect 48240 181354 48268 207674
rect 49344 183530 49372 209879
rect 49422 208090 49478 208099
rect 49422 208025 49478 208034
rect 49332 183524 49384 183530
rect 49332 183466 49384 183472
rect 49436 181490 49464 208025
rect 49528 195974 49556 228153
rect 49620 208371 49648 286282
rect 111708 286068 111760 286074
rect 111708 286010 111760 286016
rect 108948 286000 109000 286006
rect 108946 285968 108948 285977
rect 111720 285977 111748 286010
rect 109000 285968 109002 285977
rect 104808 285932 104860 285938
rect 108946 285903 109002 285912
rect 111706 285968 111762 285977
rect 111706 285903 111762 285912
rect 104808 285874 104860 285880
rect 86868 285864 86920 285870
rect 86868 285806 86920 285812
rect 81348 285796 81400 285802
rect 81348 285738 81400 285744
rect 79968 285728 80020 285734
rect 79966 285696 79968 285705
rect 81360 285705 81388 285738
rect 86880 285705 86908 285806
rect 104820 285705 104848 285874
rect 121380 285705 121408 286418
rect 136548 286408 136600 286414
rect 136546 286376 136548 286385
rect 136600 286376 136602 286385
rect 136546 286311 136602 286320
rect 133788 286272 133840 286278
rect 133788 286214 133840 286220
rect 132316 286204 132368 286210
rect 132316 286146 132368 286152
rect 126888 286136 126940 286142
rect 126886 286104 126888 286113
rect 132328 286113 132356 286146
rect 133800 286113 133828 286214
rect 126940 286104 126942 286113
rect 126886 286039 126942 286048
rect 132314 286104 132370 286113
rect 132314 286039 132370 286048
rect 133786 286104 133842 286113
rect 133786 286039 133842 286048
rect 80020 285696 80022 285705
rect 79966 285631 80022 285640
rect 81346 285696 81402 285705
rect 81346 285631 81402 285640
rect 86866 285696 86922 285705
rect 86866 285631 86922 285640
rect 89626 285696 89682 285705
rect 89626 285631 89682 285640
rect 93674 285696 93730 285705
rect 93674 285631 93730 285640
rect 102046 285696 102102 285705
rect 102046 285631 102102 285640
rect 104806 285696 104862 285705
rect 104806 285631 104862 285640
rect 106186 285696 106242 285705
rect 121366 285696 121422 285705
rect 106186 285631 106242 285640
rect 113824 285660 113876 285666
rect 89640 285326 89668 285631
rect 93688 285394 93716 285631
rect 102060 285530 102088 285631
rect 106200 285598 106228 285631
rect 121366 285631 121422 285640
rect 113824 285602 113876 285608
rect 106188 285592 106240 285598
rect 106188 285534 106240 285540
rect 102048 285524 102100 285530
rect 102048 285466 102100 285472
rect 96160 285456 96212 285462
rect 96160 285398 96212 285404
rect 93676 285388 93728 285394
rect 93676 285330 93728 285336
rect 89628 285320 89680 285326
rect 89628 285262 89680 285268
rect 96172 285161 96200 285398
rect 113836 285161 113864 285602
rect 128728 285252 128780 285258
rect 128728 285194 128780 285200
rect 123576 285184 123628 285190
rect 96158 285152 96214 285161
rect 96158 285087 96214 285096
rect 113822 285152 113878 285161
rect 123574 285152 123576 285161
rect 128740 285161 128768 285194
rect 123628 285152 123630 285161
rect 113822 285087 113878 285096
rect 118608 285116 118660 285122
rect 123574 285087 123630 285096
rect 128726 285152 128782 285161
rect 128726 285087 128782 285096
rect 118608 285058 118660 285064
rect 98552 285048 98604 285054
rect 98550 285016 98552 285025
rect 118620 285025 118648 285058
rect 98604 285016 98606 285025
rect 91192 284980 91244 284986
rect 98550 284951 98606 284960
rect 118606 285016 118662 285025
rect 118606 284951 118662 284960
rect 91192 284922 91244 284928
rect 91204 284889 91232 284922
rect 91190 284880 91246 284889
rect 91190 284815 91246 284824
rect 137296 283626 137324 286418
rect 139320 285705 139348 288390
rect 142080 285705 142108 291178
rect 144840 285705 144868 293966
rect 146220 285705 146248 296686
rect 148980 285705 149008 300834
rect 151740 285705 151768 303622
rect 154488 290488 154540 290494
rect 154488 290430 154540 290436
rect 154500 285705 154528 290430
rect 157260 285705 157288 309130
rect 169760 286544 169812 286550
rect 169760 286486 169812 286492
rect 170680 286544 170732 286550
rect 170680 286486 170732 286492
rect 169668 286476 169720 286482
rect 169668 286418 169720 286424
rect 169680 286249 169708 286418
rect 169666 286240 169722 286249
rect 169666 286175 169722 286184
rect 139306 285696 139362 285705
rect 139306 285631 139362 285640
rect 142066 285696 142122 285705
rect 142066 285631 142122 285640
rect 144826 285696 144882 285705
rect 144826 285631 144882 285640
rect 146206 285696 146262 285705
rect 146206 285631 146262 285640
rect 148966 285696 149022 285705
rect 148966 285631 149022 285640
rect 151726 285696 151782 285705
rect 151726 285631 151782 285640
rect 154486 285696 154542 285705
rect 154486 285631 154542 285640
rect 157246 285696 157302 285705
rect 157246 285631 157302 285640
rect 169772 284918 169800 286486
rect 170692 286385 170720 286486
rect 170678 286376 170734 286385
rect 180720 286346 180748 377295
rect 188448 377262 188476 458186
rect 188528 447160 188580 447166
rect 188528 447102 188580 447108
rect 188540 377330 188568 447102
rect 188632 444378 188660 464102
rect 189078 459232 189134 459241
rect 189078 459167 189134 459176
rect 189092 458318 189120 459167
rect 189080 458312 189132 458318
rect 189080 458254 189132 458260
rect 188620 444372 188672 444378
rect 188620 444314 188672 444320
rect 188620 441652 188672 441658
rect 188620 441594 188672 441600
rect 188632 377398 188660 441594
rect 188712 437504 188764 437510
rect 188712 437446 188764 437452
rect 188724 377534 188752 437446
rect 188804 431996 188856 432002
rect 188804 431938 188856 431944
rect 188816 377602 188844 431938
rect 188896 426488 188948 426494
rect 188896 426430 188948 426436
rect 188908 378622 188936 426430
rect 188988 422340 189040 422346
rect 188988 422282 189040 422288
rect 188896 378616 188948 378622
rect 188896 378558 188948 378564
rect 189000 377670 189028 422282
rect 189078 399392 189134 399401
rect 189078 399327 189134 399336
rect 189092 398886 189120 399327
rect 189080 398880 189132 398886
rect 189080 398822 189132 398828
rect 189078 397760 189134 397769
rect 189078 397695 189134 397704
rect 189092 397526 189120 397695
rect 189080 397520 189132 397526
rect 189080 397462 189132 397468
rect 189078 396400 189134 396409
rect 189078 396335 189134 396344
rect 189092 396234 189120 396335
rect 189080 396228 189132 396234
rect 189080 396170 189132 396176
rect 189446 394904 189502 394913
rect 189446 394839 189502 394848
rect 189460 394738 189488 394839
rect 189448 394732 189500 394738
rect 189448 394674 189500 394680
rect 189078 393680 189134 393689
rect 189078 393615 189134 393624
rect 189092 393378 189120 393615
rect 189080 393372 189132 393378
rect 189080 393314 189132 393320
rect 188988 377664 189040 377670
rect 188988 377606 189040 377612
rect 188804 377596 188856 377602
rect 188804 377538 188856 377544
rect 188712 377528 188764 377534
rect 188712 377470 188764 377476
rect 188620 377392 188672 377398
rect 188620 377334 188672 377340
rect 188528 377324 188580 377330
rect 188528 377266 188580 377272
rect 188436 377256 188488 377262
rect 188436 377198 188488 377204
rect 170678 286311 170734 286320
rect 180708 286340 180760 286346
rect 180708 286282 180760 286288
rect 169760 284912 169812 284918
rect 169760 284854 169812 284860
rect 180720 284073 180748 286282
rect 186688 286272 186740 286278
rect 186688 286214 186740 286220
rect 180706 284064 180762 284073
rect 180706 283999 180762 284008
rect 137284 283620 137336 283626
rect 137284 283562 137336 283568
rect 186700 282878 186728 286214
rect 186780 286204 186832 286210
rect 186780 286146 186832 286152
rect 186688 282872 186740 282878
rect 186688 282814 186740 282820
rect 186792 280158 186820 286146
rect 186964 286136 187016 286142
rect 186964 286078 187016 286084
rect 186780 280152 186832 280158
rect 186780 280094 186832 280100
rect 186976 274650 187004 286078
rect 188804 286000 188856 286006
rect 188804 285942 188856 285948
rect 187332 285932 187384 285938
rect 187332 285874 187384 285880
rect 186964 274644 187016 274650
rect 186964 274586 187016 274592
rect 186964 271924 187016 271930
rect 186964 271866 187016 271872
rect 186976 209774 187004 271866
rect 187056 259480 187108 259486
rect 187056 259422 187108 259428
rect 186884 209746 187004 209774
rect 49606 208362 49662 208371
rect 49606 208297 49662 208306
rect 49620 207738 49648 208297
rect 49608 207732 49660 207738
rect 49608 207674 49660 207680
rect 128360 199572 128412 199578
rect 128360 199514 128412 199520
rect 120080 199504 120132 199510
rect 70582 199472 70638 199481
rect 70582 199407 70638 199416
rect 77758 199472 77814 199481
rect 77758 199407 77814 199416
rect 78862 199472 78918 199481
rect 78862 199407 78918 199416
rect 88614 199472 88670 199481
rect 88614 199407 88670 199416
rect 91190 199472 91246 199481
rect 91190 199407 91246 199416
rect 103702 199472 103758 199481
rect 111062 199472 111118 199481
rect 103702 199407 103758 199416
rect 110420 199436 110472 199442
rect 70596 199034 70624 199407
rect 77772 199102 77800 199407
rect 78876 199170 78904 199407
rect 88628 199238 88656 199407
rect 91204 199306 91232 199407
rect 91192 199300 91244 199306
rect 91192 199242 91244 199248
rect 88616 199232 88668 199238
rect 88616 199174 88668 199180
rect 78864 199164 78916 199170
rect 78864 199106 78916 199112
rect 77760 199096 77812 199102
rect 77760 199038 77812 199044
rect 70584 199028 70636 199034
rect 70584 198970 70636 198976
rect 103716 198966 103744 199407
rect 120080 199446 120132 199452
rect 111062 199407 111118 199416
rect 110420 199378 110472 199384
rect 103704 198960 103756 198966
rect 103704 198902 103756 198908
rect 82544 198892 82596 198898
rect 82544 198834 82596 198840
rect 80152 198824 80204 198830
rect 80152 198766 80204 198772
rect 80164 198665 80192 198766
rect 81348 198756 81400 198762
rect 81348 198698 81400 198704
rect 81360 198665 81388 198698
rect 82556 198665 82584 198834
rect 110432 198694 110460 199378
rect 111076 199374 111104 199407
rect 111064 199368 111116 199374
rect 111064 199310 111116 199316
rect 86224 198688 86276 198694
rect 71870 198656 71926 198665
rect 71870 198591 71926 198600
rect 75550 198656 75606 198665
rect 75550 198591 75606 198600
rect 76838 198656 76894 198665
rect 76838 198591 76894 198600
rect 80150 198656 80206 198665
rect 80150 198591 80206 198600
rect 81346 198656 81402 198665
rect 81346 198591 81402 198600
rect 82542 198656 82598 198665
rect 82542 198591 82598 198600
rect 84566 198656 84622 198665
rect 84566 198591 84622 198600
rect 86222 198656 86224 198665
rect 110420 198688 110472 198694
rect 86276 198656 86278 198665
rect 86222 198591 86278 198600
rect 87970 198656 88026 198665
rect 87970 198591 88026 198600
rect 92846 198656 92902 198665
rect 92846 198591 92902 198600
rect 93582 198656 93638 198665
rect 93582 198591 93638 198600
rect 95974 198656 96030 198665
rect 95974 198591 96030 198600
rect 104438 198656 104494 198665
rect 104438 198591 104494 198600
rect 105910 198656 105966 198665
rect 105910 198591 105912 198600
rect 71884 198490 71912 198591
rect 71872 198484 71924 198490
rect 71872 198426 71924 198432
rect 73434 198384 73490 198393
rect 73434 198319 73490 198328
rect 67546 198248 67602 198257
rect 67546 198183 67602 198192
rect 66166 197432 66222 197441
rect 66166 197367 66222 197376
rect 49516 195968 49568 195974
rect 49516 195910 49568 195916
rect 66180 183462 66208 197367
rect 67560 190466 67588 198183
rect 69662 197976 69718 197985
rect 69662 197911 69718 197920
rect 68926 197432 68982 197441
rect 68926 197367 68982 197376
rect 67548 190460 67600 190466
rect 67548 190402 67600 190408
rect 68940 189038 68968 197367
rect 69676 195906 69704 197911
rect 73448 196654 73476 198319
rect 74354 198248 74410 198257
rect 74354 198183 74410 198192
rect 73436 196648 73488 196654
rect 73436 196590 73488 196596
rect 69664 195900 69716 195906
rect 69664 195842 69716 195848
rect 74368 191826 74396 198183
rect 75564 198014 75592 198591
rect 75552 198008 75604 198014
rect 75552 197950 75604 197956
rect 76852 197878 76880 198591
rect 83646 198248 83702 198257
rect 83646 198183 83702 198192
rect 76840 197872 76892 197878
rect 76840 197814 76892 197820
rect 78586 197432 78642 197441
rect 78586 197367 78642 197376
rect 81254 197432 81310 197441
rect 81254 197367 81310 197376
rect 74356 191820 74408 191826
rect 74356 191762 74408 191768
rect 68928 189032 68980 189038
rect 68928 188974 68980 188980
rect 78600 187678 78628 197367
rect 81268 193186 81296 197367
rect 83660 196518 83688 198183
rect 84580 197130 84608 198591
rect 85854 198520 85910 198529
rect 85854 198455 85910 198464
rect 85868 197198 85896 198455
rect 85856 197192 85908 197198
rect 85856 197134 85908 197140
rect 84568 197124 84620 197130
rect 84568 197066 84620 197072
rect 87984 197062 88012 198591
rect 88246 198520 88302 198529
rect 88246 198455 88302 198464
rect 89534 198520 89590 198529
rect 89534 198455 89590 198464
rect 90822 198520 90878 198529
rect 90822 198455 90878 198464
rect 87972 197056 88024 197062
rect 87972 196998 88024 197004
rect 88260 196858 88288 198455
rect 89548 196994 89576 198455
rect 89536 196988 89588 196994
rect 89536 196930 89588 196936
rect 90836 196926 90864 198455
rect 92860 198422 92888 198591
rect 92848 198416 92900 198422
rect 92848 198358 92900 198364
rect 93596 198354 93624 198591
rect 93584 198348 93636 198354
rect 93584 198290 93636 198296
rect 95988 198286 96016 198591
rect 98366 198520 98422 198529
rect 98366 198455 98422 198464
rect 100022 198520 100078 198529
rect 100022 198455 100078 198464
rect 100942 198520 100998 198529
rect 100942 198455 100998 198464
rect 102230 198520 102286 198529
rect 102230 198455 102286 198464
rect 103334 198520 103390 198529
rect 103334 198455 103390 198464
rect 95976 198280 96028 198286
rect 95976 198222 96028 198228
rect 98380 198218 98408 198455
rect 98368 198212 98420 198218
rect 98368 198154 98420 198160
rect 90824 196920 90876 196926
rect 100036 196897 100064 198455
rect 100956 198150 100984 198455
rect 100944 198144 100996 198150
rect 100944 198086 100996 198092
rect 90824 196862 90876 196868
rect 100022 196888 100078 196897
rect 88248 196852 88300 196858
rect 100022 196823 100078 196832
rect 88248 196794 88300 196800
rect 102244 196761 102272 198455
rect 103348 197033 103376 198455
rect 103334 197024 103390 197033
rect 103334 196959 103390 196968
rect 102230 196752 102286 196761
rect 102230 196687 102286 196696
rect 104452 196625 104480 198591
rect 105964 198591 105966 198600
rect 106094 198656 106150 198665
rect 106094 198591 106150 198600
rect 108486 198656 108542 198665
rect 110420 198630 110472 198636
rect 113638 198656 113694 198665
rect 108486 198591 108542 198600
rect 113638 198591 113694 198600
rect 117042 198656 117098 198665
rect 117042 198591 117098 198600
rect 118422 198656 118478 198665
rect 118422 198591 118478 198600
rect 105912 198562 105964 198568
rect 106108 198082 106136 198591
rect 108500 198558 108528 198591
rect 108488 198552 108540 198558
rect 108488 198494 108540 198500
rect 106096 198076 106148 198082
rect 106096 198018 106148 198024
rect 107014 197976 107070 197985
rect 107014 197911 107070 197920
rect 108578 197976 108634 197985
rect 108578 197911 108634 197920
rect 109222 197976 109278 197985
rect 113652 197946 113680 198591
rect 109222 197911 109278 197920
rect 113640 197940 113692 197946
rect 104438 196616 104494 196625
rect 104438 196551 104494 196560
rect 83648 196512 83700 196518
rect 83648 196454 83700 196460
rect 107028 195838 107056 197911
rect 107016 195832 107068 195838
rect 107016 195774 107068 195780
rect 108592 195770 108620 197911
rect 108580 195764 108632 195770
rect 108580 195706 108632 195712
rect 109236 195702 109264 197911
rect 113640 197882 113692 197888
rect 117056 196722 117084 198591
rect 118436 196790 118464 198591
rect 120092 197878 120120 199446
rect 128372 198694 128400 199514
rect 121000 198688 121052 198694
rect 120998 198656 121000 198665
rect 128360 198688 128412 198694
rect 121052 198656 121054 198665
rect 120998 198591 121054 198600
rect 123574 198656 123630 198665
rect 123574 198591 123630 198600
rect 126610 198656 126666 198665
rect 128360 198630 128412 198636
rect 128910 198656 128966 198665
rect 126610 198591 126666 198600
rect 128910 198591 128966 198600
rect 146022 198656 146078 198665
rect 146022 198591 146078 198600
rect 153382 198656 153438 198665
rect 153382 198591 153438 198600
rect 173438 198656 173494 198665
rect 173438 198591 173494 198600
rect 123588 197878 123616 198591
rect 120080 197872 120132 197878
rect 120080 197814 120132 197820
rect 123576 197872 123628 197878
rect 123576 197814 123628 197820
rect 118424 196784 118476 196790
rect 118424 196726 118476 196732
rect 117044 196716 117096 196722
rect 117044 196658 117096 196664
rect 126624 196586 126652 198591
rect 128924 197810 128952 198591
rect 138662 197840 138718 197849
rect 128912 197804 128964 197810
rect 138662 197775 138718 197784
rect 141238 197840 141294 197849
rect 141238 197775 141294 197784
rect 143446 197840 143502 197849
rect 143446 197775 143502 197784
rect 128912 197746 128964 197752
rect 133510 197704 133566 197713
rect 133510 197639 133566 197648
rect 126612 196580 126664 196586
rect 126612 196522 126664 196528
rect 109224 195696 109276 195702
rect 109224 195638 109276 195644
rect 133524 195158 133552 197639
rect 138676 195634 138704 197775
rect 138664 195628 138716 195634
rect 138664 195570 138716 195576
rect 141252 195566 141280 197775
rect 141240 195560 141292 195566
rect 141240 195502 141292 195508
rect 143460 195498 143488 197775
rect 143448 195492 143500 195498
rect 143448 195434 143500 195440
rect 146036 195430 146064 198591
rect 148598 197704 148654 197713
rect 148598 197639 148654 197648
rect 150990 197704 151046 197713
rect 150990 197639 151046 197648
rect 146024 195424 146076 195430
rect 146024 195366 146076 195372
rect 148612 195362 148640 197639
rect 148600 195356 148652 195362
rect 148600 195298 148652 195304
rect 151004 195294 151032 197639
rect 150992 195288 151044 195294
rect 150992 195230 151044 195236
rect 153396 195226 153424 198591
rect 173254 197840 173310 197849
rect 173254 197775 173310 197784
rect 155958 197432 156014 197441
rect 155958 197367 156014 197376
rect 153384 195220 153436 195226
rect 153384 195162 153436 195168
rect 133512 195152 133564 195158
rect 133512 195094 133564 195100
rect 155972 194546 156000 197367
rect 173268 196450 173296 197775
rect 173452 197334 173480 198591
rect 173440 197328 173492 197334
rect 173440 197270 173492 197276
rect 186884 196586 186912 209746
rect 186964 200796 187016 200802
rect 186964 200738 187016 200744
rect 186976 197946 187004 200738
rect 186964 197940 187016 197946
rect 186964 197882 187016 197888
rect 187068 196722 187096 259422
rect 187148 253972 187200 253978
rect 187148 253914 187200 253920
rect 187160 199374 187188 253914
rect 187240 245676 187292 245682
rect 187240 245618 187292 245624
rect 187148 199368 187200 199374
rect 187148 199310 187200 199316
rect 187252 198082 187280 245618
rect 187344 242894 187372 285874
rect 188344 285864 188396 285870
rect 188344 285806 188396 285812
rect 187332 242888 187384 242894
rect 187332 242830 187384 242836
rect 187332 213988 187384 213994
rect 187332 213930 187384 213936
rect 187344 199170 187372 213930
rect 188252 209908 188304 209914
rect 188252 209850 188304 209856
rect 187424 209840 187476 209846
rect 187424 209782 187476 209788
rect 187332 199164 187384 199170
rect 187332 199106 187384 199112
rect 187436 199102 187464 209782
rect 188160 205692 188212 205698
rect 188160 205634 188212 205640
rect 187424 199096 187476 199102
rect 187424 199038 187476 199044
rect 188172 198490 188200 205634
rect 188264 199238 188292 209850
rect 188356 206990 188384 285806
rect 188712 285592 188764 285598
rect 188712 285534 188764 285540
rect 188436 274712 188488 274718
rect 188436 274654 188488 274660
rect 188344 206984 188396 206990
rect 188344 206926 188396 206932
rect 188344 200184 188396 200190
rect 188344 200126 188396 200132
rect 188252 199232 188304 199238
rect 188252 199174 188304 199180
rect 188356 199034 188384 200126
rect 188344 199028 188396 199034
rect 188344 198970 188396 198976
rect 188160 198484 188212 198490
rect 188160 198426 188212 198432
rect 187240 198076 187292 198082
rect 187240 198018 187292 198024
rect 188448 197810 188476 274654
rect 188528 269136 188580 269142
rect 188528 269078 188580 269084
rect 188540 197878 188568 269078
rect 188620 262268 188672 262274
rect 188620 262210 188672 262216
rect 188528 197872 188580 197878
rect 188528 197814 188580 197820
rect 188436 197804 188488 197810
rect 188436 197746 188488 197752
rect 188632 196790 188660 262210
rect 188724 248402 188752 285534
rect 188816 252550 188844 285942
rect 188896 285660 188948 285666
rect 188896 285602 188948 285608
rect 188908 259418 188936 285602
rect 189078 279168 189134 279177
rect 189078 279103 189134 279112
rect 189092 278798 189120 279103
rect 189080 278792 189132 278798
rect 189080 278734 189132 278740
rect 188896 259412 188948 259418
rect 188896 259354 188948 259360
rect 188804 252544 188856 252550
rect 188804 252486 188856 252492
rect 188712 248396 188764 248402
rect 188712 248338 188764 248344
rect 188712 236020 188764 236026
rect 188712 235962 188764 235968
rect 188724 198150 188752 235962
rect 188804 230512 188856 230518
rect 188804 230454 188856 230460
rect 188816 198218 188844 230454
rect 188896 220856 188948 220862
rect 188896 220798 188948 220804
rect 188908 198354 188936 220798
rect 189078 219328 189134 219337
rect 189078 219263 189134 219272
rect 189092 218142 189120 219263
rect 189080 218136 189132 218142
rect 189080 218078 189132 218084
rect 189078 217696 189134 217705
rect 189078 217631 189134 217640
rect 189092 216714 189120 217631
rect 189080 216708 189132 216714
rect 189080 216650 189132 216656
rect 189170 216336 189226 216345
rect 189170 216271 189226 216280
rect 189184 215422 189212 216271
rect 189172 215416 189224 215422
rect 189172 215358 189224 215364
rect 188988 215348 189040 215354
rect 188988 215290 189040 215296
rect 189000 199306 189028 215290
rect 189080 213852 189132 213858
rect 189080 213794 189132 213800
rect 189092 213761 189120 213794
rect 189078 213752 189134 213761
rect 189078 213687 189134 213696
rect 189632 207052 189684 207058
rect 189632 206994 189684 207000
rect 189080 201544 189132 201550
rect 189080 201486 189132 201492
rect 188988 199300 189040 199306
rect 188988 199242 189040 199248
rect 188896 198348 188948 198354
rect 188896 198290 188948 198296
rect 188804 198212 188856 198218
rect 188804 198154 188856 198160
rect 188712 198144 188764 198150
rect 188712 198086 188764 198092
rect 189092 197305 189120 201486
rect 189644 199617 189672 206994
rect 189630 199608 189686 199617
rect 189630 199543 189686 199552
rect 189078 197296 189134 197305
rect 189078 197231 189134 197240
rect 188620 196784 188672 196790
rect 188620 196726 188672 196732
rect 187056 196716 187108 196722
rect 187056 196658 187108 196664
rect 186872 196580 186924 196586
rect 186872 196522 186924 196528
rect 173256 196444 173308 196450
rect 173256 196386 173308 196392
rect 155960 194540 156012 194546
rect 155960 194482 156012 194488
rect 81256 193180 81308 193186
rect 81256 193122 81308 193128
rect 78588 187672 78640 187678
rect 78588 187614 78640 187620
rect 66168 183456 66220 183462
rect 66168 183398 66220 183404
rect 49424 181484 49476 181490
rect 49424 181426 49476 181432
rect 47584 181348 47636 181354
rect 47584 181290 47636 181296
rect 48228 181348 48280 181354
rect 48228 181290 48280 181296
rect 46296 179376 46348 179382
rect 46296 179318 46348 179324
rect 46204 179240 46256 179246
rect 46204 179182 46256 179188
rect 23480 176588 23532 176594
rect 23480 176530 23532 176536
rect 3424 150408 3476 150414
rect 3424 150350 3476 150356
rect 3436 149841 3464 150350
rect 3422 149832 3478 149841
rect 3422 149767 3478 149776
rect 3240 137964 3292 137970
rect 3240 137906 3292 137912
rect 3252 136785 3280 137906
rect 3238 136776 3294 136785
rect 3238 136711 3294 136720
rect 3148 85536 3200 85542
rect 3148 85478 3200 85484
rect 3160 84697 3188 85478
rect 3146 84688 3202 84697
rect 3146 84623 3202 84632
rect 3424 45552 3476 45558
rect 3422 45520 3424 45529
rect 3476 45520 3478 45529
rect 3422 45455 3478 45464
rect 3424 6860 3476 6866
rect 3424 6802 3476 6808
rect 3436 6497 3464 6802
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 47596 3466 47624 181290
rect 48240 180878 48268 181290
rect 48228 180872 48280 180878
rect 48228 180814 48280 180820
rect 87972 180872 88024 180878
rect 87972 180814 88024 180820
rect 87984 177750 88012 180814
rect 189736 178634 189764 700334
rect 191104 565888 191156 565894
rect 191104 565830 191156 565836
rect 189814 465488 189870 465497
rect 189814 465423 189870 465432
rect 189828 336666 189856 465423
rect 189908 464976 189960 464982
rect 189908 464918 189960 464924
rect 189920 408474 189948 464918
rect 190092 464296 190144 464302
rect 190092 464238 190144 464244
rect 190000 430636 190052 430642
rect 190000 430578 190052 430584
rect 189908 408468 189960 408474
rect 189908 408410 189960 408416
rect 189908 405748 189960 405754
rect 189908 405690 189960 405696
rect 189920 378010 189948 405690
rect 190012 379001 190040 430578
rect 190104 413982 190132 464238
rect 190092 413976 190144 413982
rect 190092 413918 190144 413924
rect 190092 400240 190144 400246
rect 190092 400182 190144 400188
rect 189998 378992 190054 379001
rect 189998 378927 190054 378936
rect 190104 378078 190132 400182
rect 190184 396160 190236 396166
rect 190184 396102 190236 396108
rect 190196 379030 190224 396102
rect 190184 379024 190236 379030
rect 190184 378966 190236 378972
rect 190092 378072 190144 378078
rect 190092 378014 190144 378020
rect 189908 378004 189960 378010
rect 189908 377946 189960 377952
rect 189816 336660 189868 336666
rect 189816 336602 189868 336608
rect 189908 285320 189960 285326
rect 189908 285262 189960 285268
rect 189816 274780 189868 274786
rect 189816 274722 189868 274728
rect 189828 198937 189856 274722
rect 189920 212498 189948 285262
rect 190000 264988 190052 264994
rect 190000 264930 190052 264936
rect 189908 212492 189960 212498
rect 189908 212434 189960 212440
rect 189814 198928 189870 198937
rect 189814 198863 189870 198872
rect 190012 198422 190040 264930
rect 190092 252612 190144 252618
rect 190092 252554 190144 252560
rect 190000 198416 190052 198422
rect 190000 198358 190052 198364
rect 190104 196858 190132 252554
rect 190184 240168 190236 240174
rect 190184 240110 190236 240116
rect 190196 197130 190224 240110
rect 190276 216776 190328 216782
rect 190276 216718 190328 216724
rect 190288 197266 190316 216718
rect 190458 214840 190514 214849
rect 190458 214775 190514 214784
rect 190472 213926 190500 214775
rect 190460 213920 190512 213926
rect 190460 213862 190512 213868
rect 190368 212560 190420 212566
rect 190368 212502 190420 212508
rect 190380 199753 190408 212502
rect 190366 199744 190422 199753
rect 190366 199679 190422 199688
rect 190276 197260 190328 197266
rect 190276 197202 190328 197208
rect 190184 197124 190236 197130
rect 190184 197066 190236 197072
rect 190092 196852 190144 196858
rect 190092 196794 190144 196800
rect 191116 178974 191144 565830
rect 192484 465996 192536 466002
rect 192484 465938 192536 465944
rect 191288 465452 191340 465458
rect 191288 465394 191340 465400
rect 191196 465248 191248 465254
rect 191196 465190 191248 465196
rect 191208 358698 191236 465190
rect 191300 368490 191328 465394
rect 191288 368484 191340 368490
rect 191288 368426 191340 368432
rect 191196 358692 191248 358698
rect 191196 358634 191248 358640
rect 192496 315994 192524 465938
rect 192576 465928 192628 465934
rect 192576 465870 192628 465876
rect 192588 321502 192616 465870
rect 198188 465384 198240 465390
rect 198188 465326 198240 465332
rect 198096 465316 198148 465322
rect 198096 465258 198148 465264
rect 198004 465180 198056 465186
rect 198004 465122 198056 465128
rect 196624 464636 196676 464642
rect 196624 464578 196676 464584
rect 193864 464568 193916 464574
rect 193864 464510 193916 464516
rect 192668 464228 192720 464234
rect 192668 464170 192720 464176
rect 192680 419490 192708 464170
rect 192668 419484 192720 419490
rect 192668 419426 192720 419432
rect 192668 398880 192720 398886
rect 192668 398822 192720 398828
rect 192680 328438 192708 398822
rect 192760 397520 192812 397526
rect 192760 397462 192812 397468
rect 192772 333946 192800 397462
rect 192760 333940 192812 333946
rect 192760 333882 192812 333888
rect 193876 331226 193904 464510
rect 195244 458312 195296 458318
rect 195244 458254 195296 458260
rect 193956 426556 194008 426562
rect 193956 426498 194008 426504
rect 193968 376650 193996 426498
rect 193956 376644 194008 376650
rect 193956 376586 194008 376592
rect 193864 331220 193916 331226
rect 193864 331162 193916 331168
rect 192668 328432 192720 328438
rect 192668 328374 192720 328380
rect 192576 321496 192628 321502
rect 192576 321438 192628 321444
rect 192484 315988 192536 315994
rect 192484 315930 192536 315936
rect 195256 313206 195284 458254
rect 195336 396228 195388 396234
rect 195336 396170 195388 396176
rect 195348 340814 195376 396170
rect 195428 394732 195480 394738
rect 195428 394674 195480 394680
rect 195440 345030 195468 394674
rect 195520 393372 195572 393378
rect 195520 393314 195572 393320
rect 195532 350538 195560 393314
rect 195520 350532 195572 350538
rect 195520 350474 195572 350480
rect 195428 345024 195480 345030
rect 195428 344966 195480 344972
rect 196636 343602 196664 464578
rect 198016 353258 198044 465122
rect 198108 373998 198136 465258
rect 198200 378078 198228 465326
rect 199384 464840 199436 464846
rect 199384 464782 199436 464788
rect 198188 378072 198240 378078
rect 198188 378014 198240 378020
rect 198096 373992 198148 373998
rect 198096 373934 198148 373940
rect 199396 362846 199424 464782
rect 199384 362840 199436 362846
rect 199384 362782 199436 362788
rect 198004 353252 198056 353258
rect 198004 353194 198056 353200
rect 196624 343596 196676 343602
rect 196624 343538 196676 343544
rect 195336 340808 195388 340814
rect 195336 340750 195388 340756
rect 195244 313200 195296 313206
rect 195244 313142 195296 313148
rect 192484 286544 192536 286550
rect 192484 286486 192536 286492
rect 191380 286068 191432 286074
rect 191380 286010 191432 286016
rect 191288 285388 191340 285394
rect 191288 285330 191340 285336
rect 191196 280220 191248 280226
rect 191196 280162 191248 280168
rect 191208 199073 191236 280162
rect 191300 222154 191328 285330
rect 191392 256698 191420 286010
rect 191380 256692 191432 256698
rect 191380 256634 191432 256640
rect 191380 249824 191432 249830
rect 191380 249766 191432 249772
rect 191288 222148 191340 222154
rect 191288 222090 191340 222096
rect 191288 216708 191340 216714
rect 191288 216650 191340 216656
rect 191300 202842 191328 216650
rect 191288 202836 191340 202842
rect 191288 202778 191340 202784
rect 191194 199064 191250 199073
rect 191194 198999 191250 199008
rect 191392 197062 191420 249766
rect 191472 225004 191524 225010
rect 191472 224946 191524 224952
rect 191484 198286 191512 224946
rect 191564 215416 191616 215422
rect 191564 215358 191616 215364
rect 191576 209778 191604 215358
rect 191564 209772 191616 209778
rect 191564 209714 191616 209720
rect 191472 198280 191524 198286
rect 191472 198222 191524 198228
rect 191380 197056 191432 197062
rect 191380 196998 191432 197004
rect 192496 184890 192524 286486
rect 192668 286476 192720 286482
rect 192668 286418 192720 286424
rect 192576 278792 192628 278798
rect 192576 278734 192628 278740
rect 192484 184884 192536 184890
rect 192484 184826 192536 184832
rect 192588 182170 192616 278734
rect 192680 191758 192708 286418
rect 196716 285796 196768 285802
rect 196716 285738 196768 285744
rect 196624 285728 196676 285734
rect 196624 285670 196676 285676
rect 195244 285524 195296 285530
rect 195244 285466 195296 285472
rect 193956 285456 194008 285462
rect 193956 285398 194008 285404
rect 193864 259548 193916 259554
rect 193864 259490 193916 259496
rect 192760 255332 192812 255338
rect 192760 255274 192812 255280
rect 192772 196994 192800 255274
rect 192852 218136 192904 218142
rect 192852 218078 192904 218084
rect 192864 197266 192892 218078
rect 193128 218068 193180 218074
rect 193128 218010 193180 218016
rect 193140 213858 193168 218010
rect 193128 213852 193180 213858
rect 193128 213794 193180 213800
rect 192852 197260 192904 197266
rect 192852 197202 192904 197208
rect 192760 196988 192812 196994
rect 192760 196930 192812 196936
rect 193876 196926 193904 259490
rect 193968 227730 193996 285398
rect 194048 244316 194100 244322
rect 194048 244258 194100 244264
rect 193956 227724 194008 227730
rect 193956 227666 194008 227672
rect 193956 223644 194008 223650
rect 193956 223586 194008 223592
rect 193864 196920 193916 196926
rect 193864 196862 193916 196868
rect 193968 196450 193996 223586
rect 194060 197198 194088 244258
rect 195256 237386 195284 285466
rect 195244 237380 195296 237386
rect 195244 237322 195296 237328
rect 195244 227792 195296 227798
rect 195244 227734 195296 227740
rect 195256 197334 195284 227734
rect 195244 197328 195296 197334
rect 195244 197270 195296 197276
rect 194048 197192 194100 197198
rect 194048 197134 194100 197140
rect 193956 196444 194008 196450
rect 193956 196386 194008 196392
rect 192668 191752 192720 191758
rect 192668 191694 192720 191700
rect 196636 187610 196664 285670
rect 196728 194478 196756 285738
rect 196808 281580 196860 281586
rect 196808 281522 196860 281528
rect 196820 195158 196848 281522
rect 196808 195152 196860 195158
rect 196808 195094 196860 195100
rect 196716 194472 196768 194478
rect 196716 194414 196768 194420
rect 196624 187604 196676 187610
rect 196624 187546 196676 187552
rect 192576 182164 192628 182170
rect 192576 182106 192628 182112
rect 191104 178968 191156 178974
rect 191104 178910 191156 178916
rect 189724 178628 189776 178634
rect 189724 178570 189776 178576
rect 87972 177744 88024 177750
rect 201512 177721 201540 702986
rect 215944 462392 215996 462398
rect 215944 462334 215996 462340
rect 215956 377806 215984 462334
rect 215944 377800 215996 377806
rect 215944 377742 215996 377748
rect 87972 177686 88024 177692
rect 201498 177712 201554 177721
rect 201498 177647 201554 177656
rect 218072 177585 218100 703582
rect 218808 703474 218836 703582
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 218992 703474 219020 703520
rect 218808 703446 219020 703474
rect 239404 700324 239456 700330
rect 239404 700266 239456 700272
rect 262220 700324 262272 700330
rect 262220 700266 262272 700272
rect 235264 514820 235316 514826
rect 235264 514762 235316 514768
rect 235172 466472 235224 466478
rect 235172 466414 235224 466420
rect 235184 377777 235212 466414
rect 235170 377768 235226 377777
rect 235170 377703 235226 377712
rect 233884 345092 233936 345098
rect 233884 345034 233936 345040
rect 232504 309256 232556 309262
rect 232504 309198 232556 309204
rect 232516 194546 232544 309198
rect 232596 305108 232648 305114
rect 232596 305050 232648 305056
rect 232608 195226 232636 305050
rect 232688 302252 232740 302258
rect 232688 302194 232740 302200
rect 232700 195294 232728 302194
rect 232872 284368 232924 284374
rect 232872 284310 232924 284316
rect 232780 282940 232832 282946
rect 232780 282882 232832 282888
rect 232792 196897 232820 282882
rect 232884 198801 232912 284310
rect 232870 198792 232926 198801
rect 232870 198727 232926 198736
rect 232778 196888 232834 196897
rect 232778 196823 232834 196832
rect 232688 195288 232740 195294
rect 232688 195230 232740 195236
rect 232596 195220 232648 195226
rect 232596 195162 232648 195168
rect 232504 194540 232556 194546
rect 232504 194482 232556 194488
rect 233896 179042 233924 345034
rect 235172 289876 235224 289882
rect 235172 289818 235224 289824
rect 234988 285728 235040 285734
rect 234988 285670 235040 285676
rect 235000 197169 235028 285670
rect 234986 197160 235042 197169
rect 234986 197095 235042 197104
rect 235184 196761 235212 289818
rect 235170 196752 235226 196761
rect 235170 196687 235226 196696
rect 233884 179036 233936 179042
rect 233884 178978 233936 178984
rect 218058 177576 218114 177585
rect 218058 177511 218114 177520
rect 235276 175234 235304 514762
rect 239220 479596 239272 479602
rect 239220 479538 239272 479544
rect 237378 478952 237434 478961
rect 237378 478887 237380 478896
rect 237432 478887 237434 478896
rect 237380 478858 237432 478864
rect 237378 477864 237434 477873
rect 237378 477799 237434 477808
rect 237392 477562 237420 477799
rect 235540 477556 235592 477562
rect 235540 477498 235592 477504
rect 237380 477556 237432 477562
rect 237380 477498 237432 477504
rect 235354 465624 235410 465633
rect 235354 465559 235410 465568
rect 235368 325378 235396 465559
rect 235448 465112 235500 465118
rect 235448 465054 235500 465060
rect 235460 347682 235488 465054
rect 235552 376514 235580 477498
rect 237378 476776 237434 476785
rect 237378 476711 237434 476720
rect 237392 476134 237420 476711
rect 235632 476128 235684 476134
rect 235632 476070 235684 476076
rect 237380 476128 237432 476134
rect 237380 476070 237432 476076
rect 235644 379137 235672 476070
rect 237378 473784 237434 473793
rect 237378 473719 237434 473728
rect 237392 473414 237420 473719
rect 237380 473408 237432 473414
rect 237380 473350 237432 473356
rect 237470 472696 237526 472705
rect 237470 472631 237526 472640
rect 237378 472152 237434 472161
rect 235724 472116 235776 472122
rect 237484 472122 237512 472631
rect 237378 472087 237434 472096
rect 237472 472116 237524 472122
rect 235724 472058 235776 472064
rect 235630 379128 235686 379137
rect 235630 379063 235686 379072
rect 235736 376582 235764 472058
rect 237392 472054 237420 472087
rect 237472 472058 237524 472064
rect 235816 472048 235868 472054
rect 235816 471990 235868 471996
rect 237380 472048 237432 472054
rect 237380 471990 237432 471996
rect 235828 377641 235856 471990
rect 237378 469296 237434 469305
rect 237378 469231 237380 469240
rect 237432 469231 237434 469240
rect 237380 469202 237432 469208
rect 237378 467936 237434 467945
rect 235908 467900 235960 467906
rect 237378 467871 237380 467880
rect 235908 467842 235960 467848
rect 237432 467871 237434 467880
rect 237380 467842 237432 467848
rect 235920 379302 235948 467842
rect 237378 466712 237434 466721
rect 237378 466647 237434 466656
rect 237392 466478 237420 466647
rect 237380 466472 237432 466478
rect 237380 466414 237432 466420
rect 237380 465044 237432 465050
rect 237380 464986 237432 464992
rect 237392 464817 237420 464986
rect 238024 464908 238076 464914
rect 238024 464850 238076 464856
rect 237378 464808 237434 464817
rect 237378 464743 237434 464752
rect 237932 464772 237984 464778
rect 237932 464714 237984 464720
rect 237472 463004 237524 463010
rect 237472 462946 237524 462952
rect 237378 462632 237434 462641
rect 237378 462567 237434 462576
rect 237392 462398 237420 462567
rect 237380 462392 237432 462398
rect 237380 462334 237432 462340
rect 237484 459513 237512 462946
rect 237470 459504 237526 459513
rect 237470 459439 237526 459448
rect 237378 458280 237434 458289
rect 237378 458215 237380 458224
rect 237432 458215 237434 458224
rect 237380 458186 237432 458192
rect 237380 449880 237432 449886
rect 237380 449822 237432 449828
rect 237392 449585 237420 449822
rect 237378 449576 237434 449585
rect 237378 449511 237434 449520
rect 237378 447400 237434 447409
rect 237378 447335 237434 447344
rect 237392 447166 237420 447335
rect 237380 447160 237432 447166
rect 237380 447102 237432 447108
rect 237380 444372 237432 444378
rect 237380 444314 237432 444320
rect 237392 444281 237420 444314
rect 237378 444272 237434 444281
rect 237378 444207 237434 444216
rect 237378 442368 237434 442377
rect 237378 442303 237434 442312
rect 237392 441658 237420 442303
rect 237380 441652 237432 441658
rect 237380 441594 237432 441600
rect 237380 440224 237432 440230
rect 237380 440166 237432 440172
rect 237392 439521 237420 440166
rect 237378 439512 237434 439521
rect 237378 439447 237434 439456
rect 237378 437608 237434 437617
rect 237378 437543 237434 437552
rect 237392 437510 237420 437543
rect 237380 437504 237432 437510
rect 237380 437446 237432 437452
rect 237944 434353 237972 464714
rect 238036 454753 238064 464850
rect 238668 464704 238720 464710
rect 238668 464646 238720 464652
rect 238392 464500 238444 464506
rect 238392 464442 238444 464448
rect 238208 464432 238260 464438
rect 238208 464374 238260 464380
rect 238116 464364 238168 464370
rect 238116 464306 238168 464312
rect 238022 454744 238078 454753
rect 238022 454679 238078 454688
rect 238022 452704 238078 452713
rect 238022 452639 238078 452648
rect 237930 434344 237986 434353
rect 237930 434279 237986 434288
rect 237378 432168 237434 432177
rect 237378 432103 237434 432112
rect 237392 432002 237420 432103
rect 237380 431996 237432 432002
rect 237380 431938 237432 431944
rect 237378 431216 237434 431225
rect 237378 431151 237434 431160
rect 237392 430642 237420 431151
rect 237380 430636 237432 430642
rect 237380 430578 237432 430584
rect 237470 427136 237526 427145
rect 237470 427071 237526 427080
rect 237378 426728 237434 426737
rect 237378 426663 237434 426672
rect 237392 426562 237420 426663
rect 237380 426556 237432 426562
rect 237380 426498 237432 426504
rect 237484 426494 237512 427071
rect 237472 426488 237524 426494
rect 237472 426430 237524 426436
rect 237380 423632 237432 423638
rect 237378 423600 237380 423609
rect 237432 423600 237434 423609
rect 237378 423535 237434 423544
rect 237378 422376 237434 422385
rect 237378 422311 237380 422320
rect 237432 422311 237434 422320
rect 237380 422282 237432 422288
rect 237380 419484 237432 419490
rect 237380 419426 237432 419432
rect 237392 419257 237420 419426
rect 237378 419248 237434 419257
rect 237378 419183 237434 419192
rect 237378 416936 237434 416945
rect 237378 416871 237434 416880
rect 237392 416838 237420 416871
rect 237380 416832 237432 416838
rect 237380 416774 237432 416780
rect 237378 415984 237434 415993
rect 237378 415919 237434 415928
rect 237392 415478 237420 415919
rect 237380 415472 237432 415478
rect 237380 415414 237432 415420
rect 237380 413976 237432 413982
rect 237378 413944 237380 413953
rect 237432 413944 237434 413953
rect 237378 413879 237434 413888
rect 237378 411904 237434 411913
rect 237378 411839 237434 411848
rect 237392 411330 237420 411839
rect 237930 411360 237986 411369
rect 237380 411324 237432 411330
rect 237930 411295 237986 411304
rect 237380 411266 237432 411272
rect 237378 408504 237434 408513
rect 237378 408439 237380 408448
rect 237432 408439 237434 408448
rect 237380 408410 237432 408416
rect 237838 407144 237894 407153
rect 237838 407079 237894 407088
rect 237378 405784 237434 405793
rect 237378 405719 237380 405728
rect 237432 405719 237434 405728
rect 237380 405690 237432 405696
rect 237378 401840 237434 401849
rect 237378 401775 237434 401784
rect 237392 401674 237420 401775
rect 237380 401668 237432 401674
rect 237380 401610 237432 401616
rect 237378 400752 237434 400761
rect 237378 400687 237434 400696
rect 237392 400246 237420 400687
rect 237380 400240 237432 400246
rect 237380 400182 237432 400188
rect 237470 396672 237526 396681
rect 237470 396607 237526 396616
rect 237378 396264 237434 396273
rect 237378 396199 237434 396208
rect 237392 396166 237420 396199
rect 237380 396160 237432 396166
rect 237380 396102 237432 396108
rect 237484 396098 237512 396607
rect 237472 396092 237524 396098
rect 237472 396034 237524 396040
rect 237378 392184 237434 392193
rect 237378 392119 237434 392128
rect 237392 392018 237420 392119
rect 237380 392012 237432 392018
rect 237380 391954 237432 391960
rect 237378 390688 237434 390697
rect 237378 390623 237434 390632
rect 237392 390590 237420 390623
rect 237380 390584 237432 390590
rect 237380 390526 237432 390532
rect 237380 389156 237432 389162
rect 237380 389098 237432 389104
rect 237392 388793 237420 389098
rect 237378 388784 237434 388793
rect 237378 388719 237434 388728
rect 237378 386608 237434 386617
rect 237378 386543 237434 386552
rect 237392 386442 237420 386543
rect 237380 386436 237432 386442
rect 237380 386378 237432 386384
rect 237378 385520 237434 385529
rect 237378 385455 237434 385464
rect 237392 385082 237420 385455
rect 237380 385076 237432 385082
rect 237380 385018 237432 385024
rect 237380 383648 237432 383654
rect 237378 383616 237380 383625
rect 237432 383616 237434 383625
rect 237378 383551 237434 383560
rect 237470 381576 237526 381585
rect 237470 381511 237526 381520
rect 237378 381032 237434 381041
rect 237378 380967 237434 380976
rect 237392 380934 237420 380967
rect 237380 380928 237432 380934
rect 237380 380870 237432 380876
rect 235908 379296 235960 379302
rect 235908 379238 235960 379244
rect 237484 378894 237512 381511
rect 237472 378888 237524 378894
rect 237472 378830 237524 378836
rect 237852 378826 237880 407079
rect 237944 380186 237972 411295
rect 237932 380180 237984 380186
rect 237932 380122 237984 380128
rect 238036 379234 238064 452639
rect 238128 393961 238156 464306
rect 238220 398857 238248 464374
rect 238298 446448 238354 446457
rect 238298 446383 238354 446392
rect 238206 398848 238262 398857
rect 238206 398783 238262 398792
rect 238114 393952 238170 393961
rect 238114 393887 238170 393896
rect 238024 379228 238076 379234
rect 238024 379170 238076 379176
rect 237840 378820 237892 378826
rect 237840 378762 237892 378768
rect 237380 378072 237432 378078
rect 237378 378040 237380 378049
rect 237432 378040 237434 378049
rect 237378 377975 237434 377984
rect 235814 377632 235870 377641
rect 235814 377567 235870 377576
rect 237380 377460 237432 377466
rect 237380 377402 237432 377408
rect 237392 377233 237420 377402
rect 237378 377224 237434 377233
rect 237378 377159 237434 377168
rect 238312 377097 238340 446383
rect 238404 404025 238432 464442
rect 238482 441688 238538 441697
rect 238482 441623 238538 441632
rect 238390 404016 238446 404025
rect 238390 403951 238446 403960
rect 238496 379409 238524 441623
rect 238574 436248 238630 436257
rect 238574 436183 238630 436192
rect 238482 379400 238538 379409
rect 238482 379335 238538 379344
rect 238588 377194 238616 436183
rect 238680 429185 238708 464646
rect 238666 429176 238722 429185
rect 238666 429111 238722 429120
rect 238666 421016 238722 421025
rect 238666 420951 238722 420960
rect 238680 378729 238708 420951
rect 238666 378720 238722 378729
rect 238666 378655 238722 378664
rect 238576 377188 238628 377194
rect 238576 377130 238628 377136
rect 238298 377088 238354 377097
rect 238298 377023 238354 377032
rect 237380 376712 237432 376718
rect 237378 376680 237380 376689
rect 237432 376680 237434 376689
rect 237378 376615 237434 376624
rect 235724 376576 235776 376582
rect 235724 376518 235776 376524
rect 235540 376508 235592 376514
rect 235540 376450 235592 376456
rect 238024 376032 238076 376038
rect 238024 375974 238076 375980
rect 237380 373992 237432 373998
rect 237380 373934 237432 373940
rect 237392 373697 237420 373934
rect 237378 373688 237434 373697
rect 237378 373623 237434 373632
rect 237380 372564 237432 372570
rect 237380 372506 237432 372512
rect 237392 372473 237420 372506
rect 237378 372464 237434 372473
rect 237378 372399 237434 372408
rect 237380 371204 237432 371210
rect 237380 371146 237432 371152
rect 237392 371113 237420 371146
rect 237378 371104 237434 371113
rect 237378 371039 237434 371048
rect 237380 368484 237432 368490
rect 237380 368426 237432 368432
rect 237392 368393 237420 368426
rect 237378 368384 237434 368393
rect 237378 368319 237434 368328
rect 237472 367056 237524 367062
rect 237378 367024 237434 367033
rect 237472 366998 237524 367004
rect 237378 366959 237380 366968
rect 237432 366959 237434 366968
rect 237380 366930 237432 366936
rect 237484 366489 237512 366998
rect 237470 366480 237526 366489
rect 237470 366415 237526 366424
rect 237472 362908 237524 362914
rect 237472 362850 237524 362856
rect 237380 362840 237432 362846
rect 237378 362808 237380 362817
rect 237432 362808 237434 362817
rect 237378 362743 237434 362752
rect 237484 362545 237512 362850
rect 237470 362536 237526 362545
rect 237470 362471 237526 362480
rect 237380 361548 237432 361554
rect 237380 361490 237432 361496
rect 237392 361457 237420 361490
rect 237378 361448 237434 361457
rect 237378 361383 237434 361392
rect 237380 360188 237432 360194
rect 237380 360130 237432 360136
rect 237392 360097 237420 360130
rect 237378 360088 237434 360097
rect 237378 360023 237434 360032
rect 237380 358760 237432 358766
rect 237378 358728 237380 358737
rect 237432 358728 237434 358737
rect 237378 358663 237434 358672
rect 237472 358692 237524 358698
rect 237472 358634 237524 358640
rect 237484 358465 237512 358634
rect 237470 358456 237526 358465
rect 237470 358391 237526 358400
rect 237380 357400 237432 357406
rect 237378 357368 237380 357377
rect 237432 357368 237434 357377
rect 237378 357303 237434 357312
rect 237380 356040 237432 356046
rect 237380 355982 237432 355988
rect 237392 355881 237420 355982
rect 237472 355972 237524 355978
rect 237472 355914 237524 355920
rect 237378 355872 237434 355881
rect 237378 355807 237434 355816
rect 237484 355337 237512 355914
rect 237470 355328 237526 355337
rect 237470 355263 237526 355272
rect 237380 354680 237432 354686
rect 237380 354622 237432 354628
rect 237392 354385 237420 354622
rect 237378 354376 237434 354385
rect 237378 354311 237434 354320
rect 237380 353252 237432 353258
rect 237380 353194 237432 353200
rect 237392 353025 237420 353194
rect 237378 353016 237434 353025
rect 237378 352951 237434 352960
rect 237472 351892 237524 351898
rect 237472 351834 237524 351840
rect 237380 351824 237432 351830
rect 237378 351792 237380 351801
rect 237432 351792 237434 351801
rect 237378 351727 237434 351736
rect 237484 351393 237512 351834
rect 237470 351384 237526 351393
rect 237470 351319 237526 351328
rect 237380 350532 237432 350538
rect 237380 350474 237432 350480
rect 237392 350305 237420 350474
rect 237378 350296 237434 350305
rect 237378 350231 237434 350240
rect 237380 349104 237432 349110
rect 237378 349072 237380 349081
rect 237432 349072 237434 349081
rect 237378 349007 237434 349016
rect 237380 347744 237432 347750
rect 237380 347686 237432 347692
rect 237470 347712 237526 347721
rect 235448 347676 235500 347682
rect 235448 347618 235500 347624
rect 237392 347313 237420 347686
rect 237470 347647 237472 347656
rect 237524 347647 237526 347656
rect 237472 347618 237524 347624
rect 237378 347304 237434 347313
rect 237378 347239 237434 347248
rect 237380 346384 237432 346390
rect 237380 346326 237432 346332
rect 237392 346225 237420 346326
rect 237378 346216 237434 346225
rect 237378 346151 237434 346160
rect 237380 345024 237432 345030
rect 237380 344966 237432 344972
rect 237392 344865 237420 344966
rect 237378 344856 237434 344865
rect 237378 344791 237434 344800
rect 238036 343641 238064 375974
rect 238116 365016 238168 365022
rect 238116 364958 238168 364964
rect 238022 343632 238078 343641
rect 237380 343596 237432 343602
rect 238022 343567 238078 343576
rect 237380 343538 237432 343544
rect 237392 343233 237420 343538
rect 237378 343224 237434 343233
rect 237378 343159 237434 343168
rect 237380 342236 237432 342242
rect 237380 342178 237432 342184
rect 237392 342145 237420 342178
rect 237378 342136 237434 342145
rect 237378 342071 237434 342080
rect 237380 340876 237432 340882
rect 237380 340818 237432 340824
rect 237392 340785 237420 340818
rect 237472 340808 237524 340814
rect 237378 340776 237434 340785
rect 237472 340750 237524 340756
rect 237378 340711 237434 340720
rect 237484 340241 237512 340750
rect 237470 340232 237526 340241
rect 237470 340167 237526 340176
rect 238128 339153 238156 364958
rect 238114 339144 238170 339153
rect 238114 339079 238170 339088
rect 237380 338088 237432 338094
rect 237378 338056 237380 338065
rect 237432 338056 237434 338065
rect 237378 337991 237434 338000
rect 237472 336728 237524 336734
rect 237472 336670 237524 336676
rect 237380 336660 237432 336666
rect 237380 336602 237432 336608
rect 237392 336569 237420 336602
rect 237378 336560 237434 336569
rect 237378 336495 237434 336504
rect 237484 336161 237512 336670
rect 237470 336152 237526 336161
rect 237470 336087 237526 336096
rect 237380 335300 237432 335306
rect 237380 335242 237432 335248
rect 237392 335073 237420 335242
rect 237378 335064 237434 335073
rect 237378 334999 237434 335008
rect 237380 333940 237432 333946
rect 237380 333882 237432 333888
rect 237392 333849 237420 333882
rect 237378 333840 237434 333849
rect 237378 333775 237434 333784
rect 237380 332580 237432 332586
rect 237380 332522 237432 332528
rect 237392 332489 237420 332522
rect 237472 332512 237524 332518
rect 237378 332480 237434 332489
rect 237472 332454 237524 332460
rect 237378 332415 237434 332424
rect 237484 332081 237512 332454
rect 237470 332072 237526 332081
rect 237470 332007 237526 332016
rect 237380 331220 237432 331226
rect 237380 331162 237432 331168
rect 237392 331129 237420 331162
rect 237378 331120 237434 331129
rect 237378 331055 237434 331064
rect 237472 329792 237524 329798
rect 237472 329734 237524 329740
rect 237380 329724 237432 329730
rect 237380 329666 237432 329672
rect 237392 329633 237420 329666
rect 237378 329624 237434 329633
rect 237378 329559 237434 329568
rect 237484 329089 237512 329734
rect 237470 329080 237526 329089
rect 237470 329015 237526 329024
rect 237380 328432 237432 328438
rect 237380 328374 237432 328380
rect 237392 328001 237420 328374
rect 237378 327992 237434 328001
rect 237378 327927 237434 327936
rect 237380 327072 237432 327078
rect 237378 327040 237380 327049
rect 237432 327040 237434 327049
rect 237378 326975 237434 326984
rect 237380 325644 237432 325650
rect 237380 325586 237432 325592
rect 237392 325553 237420 325586
rect 237378 325544 237434 325553
rect 237378 325479 237434 325488
rect 235356 325372 235408 325378
rect 235356 325314 235408 325320
rect 237380 325372 237432 325378
rect 237380 325314 237432 325320
rect 237392 325009 237420 325314
rect 237378 325000 237434 325009
rect 237378 324935 237434 324944
rect 237472 324964 237524 324970
rect 237472 324906 237524 324912
rect 237380 324284 237432 324290
rect 237380 324226 237432 324232
rect 237392 323921 237420 324226
rect 237378 323912 237434 323921
rect 237378 323847 237434 323856
rect 237484 322833 237512 324906
rect 237564 323604 237616 323610
rect 237564 323546 237616 323552
rect 237470 322824 237526 322833
rect 237470 322759 237526 322768
rect 237472 321564 237524 321570
rect 237472 321506 237524 321512
rect 237380 321496 237432 321502
rect 237378 321464 237380 321473
rect 237432 321464 237434 321473
rect 237378 321399 237434 321408
rect 237484 320929 237512 321506
rect 237470 320920 237526 320929
rect 237470 320855 237526 320864
rect 237380 320136 237432 320142
rect 237380 320078 237432 320084
rect 237392 319977 237420 320078
rect 237378 319968 237434 319977
rect 237378 319903 237434 319912
rect 237380 317416 237432 317422
rect 237378 317384 237380 317393
rect 237432 317384 237434 317393
rect 237378 317319 237434 317328
rect 237576 316849 237604 323546
rect 237562 316840 237618 316849
rect 237562 316775 237618 316784
rect 237380 315988 237432 315994
rect 237380 315930 237432 315936
rect 237392 315897 237420 315930
rect 237378 315888 237434 315897
rect 237378 315823 237434 315832
rect 237380 314628 237432 314634
rect 237380 314570 237432 314576
rect 237392 314537 237420 314570
rect 237378 314528 237434 314537
rect 237378 314463 237434 314472
rect 237380 313268 237432 313274
rect 237380 313210 237432 313216
rect 237392 313177 237420 313210
rect 237472 313200 237524 313206
rect 237378 313168 237434 313177
rect 237472 313142 237524 313148
rect 237378 313103 237434 313112
rect 237484 312769 237512 313142
rect 237470 312760 237526 312769
rect 237470 312695 237526 312704
rect 237380 311840 237432 311846
rect 237378 311808 237380 311817
rect 237432 311808 237434 311817
rect 237378 311743 237434 311752
rect 237378 309496 237434 309505
rect 237378 309431 237434 309440
rect 237392 309194 237420 309431
rect 237472 309256 237524 309262
rect 237470 309224 237472 309233
rect 237524 309224 237526 309233
rect 237380 309188 237432 309194
rect 237470 309159 237526 309168
rect 237380 309130 237432 309136
rect 237378 307864 237434 307873
rect 235356 307828 235408 307834
rect 237378 307799 237380 307808
rect 235356 307770 235408 307776
rect 237432 307799 237434 307808
rect 237380 307770 237432 307776
rect 235368 195702 235396 307770
rect 238022 306504 238078 306513
rect 238022 306439 238078 306448
rect 237470 305552 237526 305561
rect 237470 305487 237526 305496
rect 237484 305114 237512 305487
rect 237472 305108 237524 305114
rect 237472 305050 237524 305056
rect 235448 305040 235500 305046
rect 237380 305040 237432 305046
rect 235448 304982 235500 304988
rect 237378 305008 237380 305017
rect 237432 305008 237434 305017
rect 235460 195770 235488 304982
rect 237378 304943 237434 304952
rect 237378 303920 237434 303929
rect 237378 303855 237434 303864
rect 237392 303686 237420 303855
rect 237380 303680 237432 303686
rect 237380 303622 237432 303628
rect 237378 302424 237434 302433
rect 237378 302359 237434 302368
rect 237392 302258 237420 302359
rect 237380 302252 237432 302258
rect 237380 302194 237432 302200
rect 237470 301472 237526 301481
rect 237470 301407 237526 301416
rect 237484 300966 237512 301407
rect 235540 300960 235592 300966
rect 237472 300960 237524 300966
rect 235540 300902 235592 300908
rect 237378 300928 237434 300937
rect 235552 195838 235580 300902
rect 237472 300902 237524 300908
rect 237378 300863 237380 300872
rect 237432 300863 237434 300872
rect 237380 300834 237432 300840
rect 236734 300112 236790 300121
rect 236734 300047 236790 300056
rect 235632 298172 235684 298178
rect 235632 298114 235684 298120
rect 235644 198626 235672 298114
rect 235724 295384 235776 295390
rect 235724 295326 235776 295332
rect 235632 198620 235684 198626
rect 235632 198562 235684 198568
rect 235736 196625 235764 295326
rect 236644 292664 236696 292670
rect 236644 292606 236696 292612
rect 235908 292596 235960 292602
rect 235908 292538 235960 292544
rect 235816 227860 235868 227866
rect 235816 227802 235868 227808
rect 235828 199889 235856 227802
rect 235814 199880 235870 199889
rect 235814 199815 235870 199824
rect 235920 197033 235948 292538
rect 235906 197024 235962 197033
rect 235906 196959 235962 196968
rect 235722 196616 235778 196625
rect 235722 196551 235778 196560
rect 235540 195832 235592 195838
rect 235540 195774 235592 195780
rect 235448 195764 235500 195770
rect 235448 195706 235500 195712
rect 235356 195696 235408 195702
rect 235356 195638 235408 195644
rect 236656 179110 236684 292606
rect 236748 195362 236776 300047
rect 237378 298888 237434 298897
rect 237378 298823 237434 298832
rect 237392 298178 237420 298823
rect 237380 298172 237432 298178
rect 237380 298114 237432 298120
rect 237378 297936 237434 297945
rect 237378 297871 237434 297880
rect 236826 296984 236882 296993
rect 236826 296919 236882 296928
rect 236840 195430 236868 296919
rect 237392 296750 237420 297871
rect 237380 296744 237432 296750
rect 237380 296686 237432 296692
rect 237378 295896 237434 295905
rect 237378 295831 237434 295840
rect 237392 295390 237420 295831
rect 237380 295384 237432 295390
rect 237380 295326 237432 295332
rect 237378 294944 237434 294953
rect 237378 294879 237434 294888
rect 237392 294030 237420 294879
rect 237380 294024 237432 294030
rect 237380 293966 237432 293972
rect 236918 293856 236974 293865
rect 236918 293791 236974 293800
rect 236932 195498 236960 293791
rect 237378 292904 237434 292913
rect 237378 292839 237434 292848
rect 237392 292602 237420 292839
rect 237380 292596 237432 292602
rect 237380 292538 237432 292544
rect 237378 291816 237434 291825
rect 237378 291751 237434 291760
rect 237392 291242 237420 291751
rect 237380 291236 237432 291242
rect 237380 291178 237432 291184
rect 237010 290864 237066 290873
rect 237010 290799 237066 290808
rect 237024 195566 237052 290799
rect 238036 290494 238064 306439
rect 238024 290488 238076 290494
rect 238024 290430 238076 290436
rect 237378 289912 237434 289921
rect 237378 289847 237380 289856
rect 237432 289847 237434 289856
rect 237380 289818 237432 289824
rect 237378 288824 237434 288833
rect 237378 288759 237434 288768
rect 237392 288454 237420 288759
rect 237380 288448 237432 288454
rect 237380 288390 237432 288396
rect 237102 287736 237158 287745
rect 237102 287671 237158 287680
rect 237116 195634 237144 287671
rect 237470 286784 237526 286793
rect 237470 286719 237526 286728
rect 237380 286408 237432 286414
rect 237380 286350 237432 286356
rect 237392 285977 237420 286350
rect 237378 285968 237434 285977
rect 237378 285903 237434 285912
rect 237484 285734 237512 286719
rect 237472 285728 237524 285734
rect 237472 285670 237524 285676
rect 238668 285252 238720 285258
rect 238668 285194 238720 285200
rect 238116 285184 238168 285190
rect 238116 285126 238168 285132
rect 238024 284980 238076 284986
rect 238024 284922 238076 284928
rect 237378 284744 237434 284753
rect 237378 284679 237434 284688
rect 237392 284374 237420 284679
rect 237380 284368 237432 284374
rect 237380 284310 237432 284316
rect 237470 283792 237526 283801
rect 237470 283727 237526 283736
rect 237484 282946 237512 283727
rect 237472 282940 237524 282946
rect 237472 282882 237524 282888
rect 237380 282872 237432 282878
rect 237378 282840 237380 282849
rect 237432 282840 237434 282849
rect 237378 282775 237434 282784
rect 237378 281752 237434 281761
rect 237378 281687 237434 281696
rect 237392 281586 237420 281687
rect 237380 281580 237432 281586
rect 237380 281522 237432 281528
rect 237470 280664 237526 280673
rect 237470 280599 237526 280608
rect 237484 280226 237512 280599
rect 237472 280220 237524 280226
rect 237472 280162 237524 280168
rect 237380 280152 237432 280158
rect 237380 280094 237432 280100
rect 237392 279857 237420 280094
rect 237378 279848 237434 279857
rect 237378 279783 237434 279792
rect 237470 275632 237526 275641
rect 237470 275567 237526 275576
rect 237378 274816 237434 274825
rect 237378 274751 237380 274760
rect 237432 274751 237434 274760
rect 237380 274722 237432 274728
rect 237484 274718 237512 275567
rect 237472 274712 237524 274718
rect 237472 274654 237524 274660
rect 237380 274644 237432 274650
rect 237380 274586 237432 274592
rect 237392 273737 237420 274586
rect 237378 273728 237434 273737
rect 237378 273663 237434 273672
rect 237378 272640 237434 272649
rect 237378 272575 237434 272584
rect 237392 271930 237420 272575
rect 237380 271924 237432 271930
rect 237380 271866 237432 271872
rect 237378 269512 237434 269521
rect 237378 269447 237434 269456
rect 237392 269142 237420 269447
rect 237380 269136 237432 269142
rect 237380 269078 237432 269084
rect 237378 265568 237434 265577
rect 237378 265503 237434 265512
rect 237392 264994 237420 265503
rect 237380 264988 237432 264994
rect 237380 264930 237432 264936
rect 237378 263528 237434 263537
rect 237378 263463 237434 263472
rect 237392 262274 237420 263463
rect 237380 262268 237432 262274
rect 237380 262210 237432 262216
rect 237470 260400 237526 260409
rect 237470 260335 237526 260344
rect 237378 259584 237434 259593
rect 237378 259519 237380 259528
rect 237432 259519 237434 259528
rect 237380 259490 237432 259496
rect 237484 259486 237512 260335
rect 237472 259480 237524 259486
rect 237472 259422 237524 259428
rect 237380 259412 237432 259418
rect 237380 259354 237432 259360
rect 237392 258505 237420 259354
rect 237378 258496 237434 258505
rect 237378 258431 237434 258440
rect 237472 256692 237524 256698
rect 237472 256634 237524 256640
rect 237378 256320 237434 256329
rect 237378 256255 237434 256264
rect 237392 255338 237420 256255
rect 237484 255513 237512 256634
rect 237470 255504 237526 255513
rect 237470 255439 237526 255448
rect 237380 255332 237432 255338
rect 237380 255274 237432 255280
rect 237378 254416 237434 254425
rect 237378 254351 237434 254360
rect 237392 253978 237420 254351
rect 237380 253972 237432 253978
rect 237380 253914 237432 253920
rect 237470 253328 237526 253337
rect 237470 253263 237526 253272
rect 237484 252618 237512 253263
rect 237472 252612 237524 252618
rect 237472 252554 237524 252560
rect 237380 252544 237432 252550
rect 237378 252512 237380 252521
rect 237432 252512 237434 252521
rect 237378 252447 237434 252456
rect 237378 250336 237434 250345
rect 237378 250271 237434 250280
rect 237392 249830 237420 250271
rect 237380 249824 237432 249830
rect 237380 249766 237432 249772
rect 237380 248396 237432 248402
rect 237380 248338 237432 248344
rect 237392 247353 237420 248338
rect 237378 247344 237434 247353
rect 237378 247279 237434 247288
rect 237378 246256 237434 246265
rect 237378 246191 237434 246200
rect 237392 245682 237420 246191
rect 237380 245676 237432 245682
rect 237380 245618 237432 245624
rect 237378 245168 237434 245177
rect 237378 245103 237434 245112
rect 237392 244322 237420 245103
rect 237380 244316 237432 244322
rect 237380 244258 237432 244264
rect 237380 242888 237432 242894
rect 237380 242830 237432 242836
rect 237392 242321 237420 242830
rect 237378 242312 237434 242321
rect 237378 242247 237434 242256
rect 237378 240272 237434 240281
rect 237378 240207 237434 240216
rect 237392 240174 237420 240207
rect 237380 240168 237432 240174
rect 237380 240110 237432 240116
rect 237380 237380 237432 237386
rect 237380 237322 237432 237328
rect 237392 237289 237420 237322
rect 237378 237280 237434 237289
rect 237378 237215 237434 237224
rect 237378 236056 237434 236065
rect 237378 235991 237380 236000
rect 237432 235991 237434 236000
rect 237380 235962 237432 235968
rect 237378 231024 237434 231033
rect 237378 230959 237434 230968
rect 237392 230518 237420 230959
rect 237380 230512 237432 230518
rect 237380 230454 237432 230460
rect 237470 228984 237526 228993
rect 237470 228919 237526 228928
rect 237378 228032 237434 228041
rect 237378 227967 237434 227976
rect 237392 227866 237420 227967
rect 237380 227860 237432 227866
rect 237380 227802 237432 227808
rect 237484 227798 237512 228919
rect 237472 227792 237524 227798
rect 237472 227734 237524 227740
rect 237380 227724 237432 227730
rect 237380 227666 237432 227672
rect 237392 227089 237420 227666
rect 237378 227080 237434 227089
rect 237378 227015 237434 227024
rect 237378 225992 237434 226001
rect 237378 225927 237434 225936
rect 237392 225010 237420 225927
rect 237380 225004 237432 225010
rect 237380 224946 237432 224952
rect 237378 223952 237434 223961
rect 237378 223887 237434 223896
rect 237392 223650 237420 223887
rect 237380 223644 237432 223650
rect 237380 223586 237432 223592
rect 237930 223000 237986 223009
rect 237930 222935 237986 222944
rect 237380 222148 237432 222154
rect 237380 222090 237432 222096
rect 237392 222057 237420 222090
rect 237378 222048 237434 222057
rect 237378 221983 237434 221992
rect 237378 220960 237434 220969
rect 237378 220895 237434 220904
rect 237392 220862 237420 220895
rect 237380 220856 237432 220862
rect 237380 220798 237432 220804
rect 237378 218920 237434 218929
rect 237378 218855 237434 218864
rect 237392 218074 237420 218855
rect 237380 218068 237432 218074
rect 237380 218010 237432 218016
rect 237378 217832 237434 217841
rect 237378 217767 237434 217776
rect 237392 216782 237420 217767
rect 237380 216776 237432 216782
rect 237380 216718 237432 216724
rect 237378 215792 237434 215801
rect 237378 215727 237434 215736
rect 237392 215354 237420 215727
rect 237380 215348 237432 215354
rect 237380 215290 237432 215296
rect 237470 214840 237526 214849
rect 237470 214775 237526 214784
rect 237484 213994 237512 214775
rect 237472 213988 237524 213994
rect 237472 213930 237524 213936
rect 237380 213920 237432 213926
rect 237378 213888 237380 213897
rect 237432 213888 237434 213897
rect 237378 213823 237434 213832
rect 237378 212800 237434 212809
rect 237378 212735 237434 212744
rect 237392 212566 237420 212735
rect 237380 212560 237432 212566
rect 237380 212502 237432 212508
rect 237472 212492 237524 212498
rect 237472 212434 237524 212440
rect 237484 211993 237512 212434
rect 237470 211984 237526 211993
rect 237470 211919 237526 211928
rect 237470 210760 237526 210769
rect 237470 210695 237526 210704
rect 237484 209914 237512 210695
rect 237472 209908 237524 209914
rect 237472 209850 237524 209856
rect 237380 209840 237432 209846
rect 237378 209808 237380 209817
rect 237432 209808 237434 209817
rect 237378 209743 237434 209752
rect 237472 209772 237524 209778
rect 237472 209714 237524 209720
rect 237484 208865 237512 209714
rect 237470 208856 237526 208865
rect 237470 208791 237526 208800
rect 237378 207768 237434 207777
rect 237378 207703 237434 207712
rect 237392 207058 237420 207703
rect 237380 207052 237432 207058
rect 237380 206994 237432 207000
rect 237472 206984 237524 206990
rect 237472 206926 237524 206932
rect 237378 206680 237434 206689
rect 237378 206615 237434 206624
rect 237392 205698 237420 206615
rect 237484 205873 237512 206926
rect 237470 205864 237526 205873
rect 237470 205799 237526 205808
rect 237380 205692 237432 205698
rect 237380 205634 237432 205640
rect 237838 203688 237894 203697
rect 237838 203623 237894 203632
rect 237380 202836 237432 202842
rect 237380 202778 237432 202784
rect 237392 202745 237420 202778
rect 237378 202736 237434 202745
rect 237378 202671 237434 202680
rect 237378 201648 237434 201657
rect 237378 201583 237434 201592
rect 237392 201550 237420 201583
rect 237380 201544 237432 201550
rect 237380 201486 237432 201492
rect 237378 200696 237434 200705
rect 237378 200631 237434 200640
rect 237392 200190 237420 200631
rect 237380 200184 237432 200190
rect 237380 200126 237432 200132
rect 237852 199510 237880 203623
rect 237840 199504 237892 199510
rect 237840 199446 237892 199452
rect 237470 198656 237526 198665
rect 237470 198591 237526 198600
rect 237380 198008 237432 198014
rect 237380 197950 237432 197956
rect 237392 197713 237420 197950
rect 237378 197704 237434 197713
rect 237378 197639 237434 197648
rect 237380 197260 237432 197266
rect 237380 197202 237432 197208
rect 237392 196761 237420 197202
rect 237378 196752 237434 196761
rect 237378 196687 237434 196696
rect 237484 196518 237512 198591
rect 237944 197742 237972 222935
rect 238036 217025 238064 284922
rect 238128 270745 238156 285126
rect 238392 285116 238444 285122
rect 238392 285058 238444 285064
rect 238208 284912 238260 284918
rect 238208 284854 238260 284860
rect 238114 270736 238170 270745
rect 238114 270671 238170 270680
rect 238114 266520 238170 266529
rect 238114 266455 238170 266464
rect 238022 217016 238078 217025
rect 238022 216951 238078 216960
rect 238022 204640 238078 204649
rect 238022 204575 238078 204584
rect 238036 199442 238064 204575
rect 238128 199578 238156 266455
rect 238220 261633 238248 284854
rect 238298 278624 238354 278633
rect 238298 278559 238354 278568
rect 238206 261624 238262 261633
rect 238206 261559 238262 261568
rect 238206 257408 238262 257417
rect 238206 257343 238262 257352
rect 238220 200802 238248 257343
rect 238312 222873 238340 278559
rect 238404 264625 238432 285058
rect 238484 285048 238536 285054
rect 238484 284990 238536 284996
rect 238390 264616 238446 264625
rect 238390 264551 238446 264560
rect 238390 251288 238446 251297
rect 238390 251223 238446 251232
rect 238298 222864 238354 222873
rect 238298 222799 238354 222808
rect 238298 219872 238354 219881
rect 238298 219807 238354 219816
rect 238208 200796 238260 200802
rect 238208 200738 238260 200744
rect 238116 199572 238168 199578
rect 238116 199514 238168 199520
rect 238024 199436 238076 199442
rect 238024 199378 238076 199384
rect 238312 198830 238340 219807
rect 238300 198824 238352 198830
rect 238300 198766 238352 198772
rect 238404 198558 238432 251223
rect 238496 232257 238524 284990
rect 238576 283620 238628 283626
rect 238576 283562 238628 283568
rect 238588 267617 238616 283562
rect 238680 276865 238708 285194
rect 238666 276856 238722 276865
rect 238666 276791 238722 276800
rect 238574 267608 238630 267617
rect 238574 267543 238630 267552
rect 238574 241224 238630 241233
rect 238574 241159 238630 241168
rect 238482 232248 238538 232257
rect 238482 232183 238538 232192
rect 238482 230072 238538 230081
rect 238482 230007 238538 230016
rect 238496 198898 238524 230007
rect 238588 198966 238616 241159
rect 238666 225040 238722 225049
rect 238666 224975 238722 224984
rect 238576 198960 238628 198966
rect 238576 198902 238628 198908
rect 238484 198892 238536 198898
rect 238484 198834 238536 198840
rect 238680 198762 238708 224975
rect 238668 198756 238720 198762
rect 238668 198698 238720 198704
rect 238392 198552 238444 198558
rect 238392 198494 238444 198500
rect 237932 197736 237984 197742
rect 237932 197678 237984 197684
rect 238024 196648 238076 196654
rect 238024 196590 238076 196596
rect 237472 196512 237524 196518
rect 237472 196454 237524 196460
rect 237380 195968 237432 195974
rect 237380 195910 237432 195916
rect 237392 195673 237420 195910
rect 237472 195900 237524 195906
rect 237472 195842 237524 195848
rect 237378 195664 237434 195673
rect 237104 195628 237156 195634
rect 237378 195599 237434 195608
rect 237104 195570 237156 195576
rect 237012 195560 237064 195566
rect 237012 195502 237064 195508
rect 236920 195492 236972 195498
rect 236920 195434 236972 195440
rect 236828 195424 236880 195430
rect 236828 195366 236880 195372
rect 236736 195356 236788 195362
rect 236736 195298 236788 195304
rect 237484 194721 237512 195842
rect 237470 194712 237526 194721
rect 237470 194647 237526 194656
rect 237380 194472 237432 194478
rect 237380 194414 237432 194420
rect 237392 193633 237420 194414
rect 237378 193624 237434 193633
rect 237378 193559 237434 193568
rect 237380 193180 237432 193186
rect 237380 193122 237432 193128
rect 237392 192681 237420 193122
rect 237378 192672 237434 192681
rect 237378 192607 237434 192616
rect 237380 191820 237432 191826
rect 237380 191762 237432 191768
rect 237392 191593 237420 191762
rect 237472 191752 237524 191758
rect 237472 191694 237524 191700
rect 237378 191584 237434 191593
rect 237378 191519 237434 191528
rect 237484 190641 237512 191694
rect 237470 190632 237526 190641
rect 237470 190567 237526 190576
rect 237380 190460 237432 190466
rect 237380 190402 237432 190408
rect 237392 189689 237420 190402
rect 237378 189680 237434 189689
rect 237378 189615 237434 189624
rect 238036 185609 238064 196590
rect 238392 189032 238444 189038
rect 238392 188974 238444 188980
rect 238404 188601 238432 188974
rect 238390 188592 238446 188601
rect 238390 188527 238446 188536
rect 239128 187740 239180 187746
rect 239128 187682 239180 187688
rect 238760 187672 238812 187678
rect 238390 187640 238446 187649
rect 238760 187614 238812 187620
rect 238390 187575 238392 187584
rect 238444 187575 238446 187584
rect 238392 187546 238444 187552
rect 238772 186561 238800 187614
rect 238758 186552 238814 186561
rect 238758 186487 238814 186496
rect 238022 185600 238078 185609
rect 238022 185535 238078 185544
rect 238760 184884 238812 184890
rect 238760 184826 238812 184832
rect 238772 184521 238800 184826
rect 238758 184512 238814 184521
rect 238758 184447 238814 184456
rect 238300 183524 238352 183530
rect 238300 183466 238352 183472
rect 238312 182481 238340 183466
rect 238392 183456 238444 183462
rect 238390 183424 238392 183433
rect 238444 183424 238446 183433
rect 238390 183359 238446 183368
rect 239036 182912 239088 182918
rect 239036 182854 239088 182860
rect 238298 182472 238354 182481
rect 238298 182407 238354 182416
rect 238576 181484 238628 181490
rect 238576 181426 238628 181432
rect 238588 180577 238616 181426
rect 238574 180568 238630 180577
rect 238574 180503 238630 180512
rect 236644 179104 236696 179110
rect 236644 179046 236696 179052
rect 239048 177274 239076 182854
rect 239140 179178 239168 187682
rect 239128 179172 239180 179178
rect 239128 179114 239180 179120
rect 239232 178770 239260 479538
rect 239312 478916 239364 478922
rect 239312 478858 239364 478864
rect 239324 182782 239352 478858
rect 239312 182776 239364 182782
rect 239312 182718 239364 182724
rect 239416 182322 239444 700266
rect 262232 696946 262260 700266
rect 267660 697610 267688 703520
rect 283852 702434 283880 703520
rect 282932 702406 283880 702434
rect 278780 700392 278832 700398
rect 278780 700334 278832 700340
rect 266360 697604 266412 697610
rect 266360 697546 266412 697552
rect 267648 697604 267700 697610
rect 267648 697546 267700 697552
rect 262140 696918 262260 696946
rect 262140 694142 262168 696918
rect 259460 694136 259512 694142
rect 259460 694078 259512 694084
rect 262128 694136 262180 694142
rect 262128 694078 262180 694084
rect 259472 687290 259500 694078
rect 259380 687262 259500 687290
rect 259380 683194 259408 687262
rect 253204 683188 253256 683194
rect 253204 683130 253256 683136
rect 259368 683188 259420 683194
rect 259368 683130 259420 683136
rect 239588 656940 239640 656946
rect 239588 656882 239640 656888
rect 239496 501016 239548 501022
rect 239496 500958 239548 500964
rect 239324 182294 239444 182322
rect 239324 178809 239352 182294
rect 239404 182164 239456 182170
rect 239404 182106 239456 182112
rect 239416 181529 239444 182106
rect 239402 181520 239458 181529
rect 239402 181455 239458 181464
rect 239508 178906 239536 500958
rect 239600 179217 239628 656882
rect 253216 627910 253244 683130
rect 251824 627904 251876 627910
rect 251824 627846 251876 627852
rect 253204 627904 253256 627910
rect 253204 627846 253256 627852
rect 251836 600506 251864 627846
rect 250444 600500 250496 600506
rect 250444 600442 250496 600448
rect 251824 600500 251876 600506
rect 251824 600442 251876 600448
rect 250456 573850 250484 600442
rect 264980 579692 265032 579698
rect 264980 579634 265032 579640
rect 264992 578202 265020 579634
rect 262864 578196 262916 578202
rect 262864 578138 262916 578144
rect 264980 578196 265032 578202
rect 264980 578138 265032 578144
rect 247684 573844 247736 573850
rect 247684 573786 247736 573792
rect 250444 573844 250496 573850
rect 250444 573786 250496 573792
rect 239772 553444 239824 553450
rect 239772 553386 239824 553392
rect 239680 480956 239732 480962
rect 239680 480898 239732 480904
rect 239692 182918 239720 480898
rect 239680 182912 239732 182918
rect 239680 182854 239732 182860
rect 239680 182776 239732 182782
rect 239680 182718 239732 182724
rect 239586 179208 239642 179217
rect 239586 179143 239642 179152
rect 239496 178900 239548 178906
rect 239496 178842 239548 178848
rect 239310 178800 239366 178809
rect 239220 178764 239272 178770
rect 239310 178735 239366 178744
rect 239220 178706 239272 178712
rect 239692 178498 239720 182718
rect 239784 179353 239812 553386
rect 247696 532506 247724 573786
rect 262876 550798 262904 578138
rect 261208 550792 261260 550798
rect 261208 550734 261260 550740
rect 262864 550792 262916 550798
rect 262864 550734 262916 550740
rect 261220 548554 261248 550734
rect 259460 548548 259512 548554
rect 259460 548490 259512 548496
rect 261208 548548 261260 548554
rect 261208 548490 261260 548496
rect 259472 547874 259500 548490
rect 259380 547846 259500 547874
rect 259380 539646 259408 547846
rect 257344 539640 257396 539646
rect 257344 539582 257396 539588
rect 259368 539640 259420 539646
rect 259368 539582 259420 539588
rect 245016 532500 245068 532506
rect 245016 532442 245068 532448
rect 247684 532500 247736 532506
rect 247684 532442 247736 532448
rect 244924 523728 244976 523734
rect 244924 523670 244976 523676
rect 243636 506524 243688 506530
rect 243636 506466 243688 506472
rect 243648 504218 243676 506466
rect 242164 504212 242216 504218
rect 242164 504154 242216 504160
rect 243636 504212 243688 504218
rect 243636 504154 243688 504160
rect 240324 484084 240376 484090
rect 240324 484026 240376 484032
rect 239864 482724 239916 482730
rect 239864 482666 239916 482672
rect 239770 179344 239826 179353
rect 239770 179279 239826 179288
rect 239876 178838 239904 482666
rect 240336 478922 240364 484026
rect 240784 483812 240836 483818
rect 240784 483754 240836 483760
rect 240796 479602 240824 483754
rect 242176 482730 242204 504154
rect 244936 496874 244964 523670
rect 245028 506530 245056 532442
rect 257356 524482 257384 539582
rect 254584 524476 254636 524482
rect 254584 524418 254636 524424
rect 257344 524476 257396 524482
rect 257344 524418 257396 524424
rect 245016 506524 245068 506530
rect 245016 506466 245068 506472
rect 254596 505170 254624 524418
rect 251640 505164 251692 505170
rect 251640 505106 251692 505112
rect 254584 505164 254636 505170
rect 254584 505106 254636 505112
rect 251652 502042 251680 505106
rect 249800 502036 249852 502042
rect 249800 501978 249852 501984
rect 251640 502036 251692 502042
rect 251640 501978 251692 501984
rect 249812 497010 249840 501978
rect 247684 497004 247736 497010
rect 247684 496946 247736 496952
rect 249800 497004 249852 497010
rect 249800 496946 249852 496952
rect 242256 496868 242308 496874
rect 242256 496810 242308 496816
rect 244924 496868 244976 496874
rect 244924 496810 244976 496816
rect 242268 484090 242296 496810
rect 247696 485858 247724 496946
rect 242808 485852 242860 485858
rect 242808 485794 242860 485800
rect 247684 485852 247736 485858
rect 247684 485794 247736 485800
rect 242256 484084 242308 484090
rect 242256 484026 242308 484032
rect 242820 483818 242848 485794
rect 242808 483812 242860 483818
rect 242808 483754 242860 483760
rect 242164 482724 242216 482730
rect 242164 482666 242216 482672
rect 266372 480962 266400 697546
rect 278792 696946 278820 700334
rect 278700 696918 278820 696946
rect 278700 692850 278728 696918
rect 276756 692844 276808 692850
rect 276756 692786 276808 692792
rect 278688 692844 278740 692850
rect 278688 692786 278740 692792
rect 276768 687546 276796 692786
rect 275284 687540 275336 687546
rect 275284 687482 275336 687488
rect 276756 687540 276808 687546
rect 276756 687482 276808 687488
rect 275296 655518 275324 687482
rect 273904 655512 273956 655518
rect 273904 655454 273956 655460
rect 275284 655512 275336 655518
rect 275284 655454 275336 655460
rect 273916 638246 273944 655454
rect 272524 638240 272576 638246
rect 272524 638182 272576 638188
rect 273904 638240 273956 638246
rect 273904 638182 273956 638188
rect 272536 623830 272564 638182
rect 269764 623824 269816 623830
rect 269764 623766 269816 623772
rect 272524 623824 272576 623830
rect 272524 623766 272576 623772
rect 269776 604518 269804 623766
rect 268752 604512 268804 604518
rect 268752 604454 268804 604460
rect 269764 604512 269816 604518
rect 269764 604454 269816 604460
rect 268764 602410 268792 604454
rect 267004 602404 267056 602410
rect 267004 602346 267056 602352
rect 268752 602404 268804 602410
rect 268752 602346 268804 602352
rect 267016 579698 267044 602346
rect 282932 588470 282960 702406
rect 332520 700330 332548 703520
rect 348804 700398 348832 703520
rect 348792 700392 348844 700398
rect 348792 700334 348844 700340
rect 332508 700324 332560 700330
rect 332508 700266 332560 700272
rect 397472 699990 397500 703520
rect 413664 700534 413692 703520
rect 413652 700528 413704 700534
rect 413652 700470 413704 700476
rect 420920 700528 420972 700534
rect 420920 700470 420972 700476
rect 397460 699984 397512 699990
rect 397460 699926 397512 699932
rect 399300 699984 399352 699990
rect 399300 699926 399352 699932
rect 399312 695502 399340 699926
rect 399300 695496 399352 695502
rect 399300 695438 399352 695444
rect 400956 695496 401008 695502
rect 400956 695438 401008 695444
rect 400968 691150 400996 695438
rect 420932 694210 420960 700470
rect 420920 694204 420972 694210
rect 420920 694146 420972 694152
rect 424324 694204 424376 694210
rect 424324 694146 424376 694152
rect 400956 691144 401008 691150
rect 400956 691086 401008 691092
rect 401968 691144 402020 691150
rect 401968 691086 402020 691092
rect 401980 684554 402008 691086
rect 424336 685166 424364 694146
rect 462332 690742 462360 703520
rect 478524 702434 478552 703520
rect 477512 702406 478552 702434
rect 477512 694822 477540 702406
rect 527192 700330 527220 703520
rect 543476 702434 543504 703520
rect 542372 702406 543504 702434
rect 527180 700324 527232 700330
rect 527180 700266 527232 700272
rect 538220 700324 538272 700330
rect 538220 700266 538272 700272
rect 477500 694816 477552 694822
rect 477500 694758 477552 694764
rect 480260 694816 480312 694822
rect 480260 694758 480312 694764
rect 462320 690736 462372 690742
rect 462320 690678 462372 690684
rect 465172 690736 465224 690742
rect 465172 690678 465224 690684
rect 465184 688226 465212 690678
rect 465172 688220 465224 688226
rect 465172 688162 465224 688168
rect 471244 688220 471296 688226
rect 471244 688162 471296 688168
rect 424324 685160 424376 685166
rect 424324 685102 424376 685108
rect 447784 685160 447836 685166
rect 447784 685102 447836 685108
rect 401968 684548 402020 684554
rect 401968 684490 402020 684496
rect 405004 684480 405056 684486
rect 405004 684422 405056 684428
rect 405016 626550 405044 684422
rect 447796 664494 447824 685102
rect 471256 681426 471284 688162
rect 480272 687954 480300 694758
rect 480260 687948 480312 687954
rect 480260 687890 480312 687896
rect 490564 687948 490616 687954
rect 490564 687890 490616 687896
rect 471244 681420 471296 681426
rect 471244 681362 471296 681368
rect 474648 681420 474700 681426
rect 474648 681362 474700 681368
rect 474660 677550 474688 681362
rect 474648 677544 474700 677550
rect 474648 677486 474700 677492
rect 478144 677544 478196 677550
rect 478144 677486 478196 677492
rect 478156 672790 478184 677486
rect 478144 672784 478196 672790
rect 478144 672726 478196 672732
rect 483664 672784 483716 672790
rect 483664 672726 483716 672732
rect 483676 664494 483704 672726
rect 490576 665174 490604 687890
rect 490564 665168 490616 665174
rect 490564 665110 490616 665116
rect 493324 665168 493376 665174
rect 493324 665110 493376 665116
rect 447784 664488 447836 664494
rect 447784 664430 447836 664436
rect 460204 664488 460256 664494
rect 460204 664430 460256 664436
rect 483664 664488 483716 664494
rect 483664 664430 483716 664436
rect 460216 656334 460244 664430
rect 460204 656328 460256 656334
rect 460204 656270 460256 656276
rect 462320 656328 462372 656334
rect 462320 656270 462372 656276
rect 462332 653206 462360 656270
rect 462320 653200 462372 653206
rect 462320 653142 462372 653148
rect 465448 653200 465500 653206
rect 465448 653142 465500 653148
rect 465460 650690 465488 653142
rect 465448 650684 465500 650690
rect 465448 650626 465500 650632
rect 480904 650684 480956 650690
rect 480904 650626 480956 650632
rect 480916 641102 480944 650626
rect 480904 641096 480956 641102
rect 480904 641038 480956 641044
rect 493336 641034 493364 665110
rect 497464 664488 497516 664494
rect 497464 664430 497516 664436
rect 497476 654838 497504 664430
rect 497464 654832 497516 654838
rect 497464 654774 497516 654780
rect 508504 654832 508556 654838
rect 508504 654774 508556 654780
rect 494704 641096 494756 641102
rect 494704 641038 494756 641044
rect 493324 641028 493376 641034
rect 493324 640970 493376 640976
rect 494716 636886 494744 641038
rect 507124 641028 507176 641034
rect 507124 640970 507176 640976
rect 494704 636880 494756 636886
rect 494704 636822 494756 636828
rect 505744 636880 505796 636886
rect 505744 636822 505796 636828
rect 405004 626544 405056 626550
rect 405004 626486 405056 626492
rect 407764 626544 407816 626550
rect 407764 626486 407816 626492
rect 407776 613086 407804 626486
rect 505756 623082 505784 636822
rect 505744 623076 505796 623082
rect 505744 623018 505796 623024
rect 407764 613080 407816 613086
rect 407764 613022 407816 613028
rect 409236 613080 409288 613086
rect 409236 613022 409288 613028
rect 409248 609958 409276 613022
rect 409236 609952 409288 609958
rect 409236 609894 409288 609900
rect 410524 609952 410576 609958
rect 410524 609894 410576 609900
rect 410536 600302 410564 609894
rect 507136 607918 507164 640970
rect 508516 633758 508544 654774
rect 508504 633752 508556 633758
rect 508504 633694 508556 633700
rect 511264 633752 511316 633758
rect 511264 633694 511316 633700
rect 511276 624442 511304 633694
rect 511264 624436 511316 624442
rect 511264 624378 511316 624384
rect 521660 624436 521712 624442
rect 521660 624378 521712 624384
rect 521672 616826 521700 624378
rect 522304 623076 522356 623082
rect 522304 623018 522356 623024
rect 521660 616820 521712 616826
rect 521660 616762 521712 616768
rect 522316 614242 522344 623018
rect 525156 616820 525208 616826
rect 525156 616762 525208 616768
rect 522304 614236 522356 614242
rect 522304 614178 522356 614184
rect 525064 614236 525116 614242
rect 525064 614178 525116 614184
rect 507124 607912 507176 607918
rect 507124 607854 507176 607860
rect 518900 607912 518952 607918
rect 518900 607854 518952 607860
rect 518912 603158 518940 607854
rect 518900 603152 518952 603158
rect 518900 603094 518952 603100
rect 522856 603152 522908 603158
rect 522856 603094 522908 603100
rect 410524 600296 410576 600302
rect 410524 600238 410576 600244
rect 411904 600296 411956 600302
rect 411904 600238 411956 600244
rect 411916 595134 411944 600238
rect 522868 596873 522896 603094
rect 522854 596864 522910 596873
rect 522854 596799 522910 596808
rect 411904 595128 411956 595134
rect 411904 595070 411956 595076
rect 414664 595128 414716 595134
rect 414664 595070 414716 595076
rect 282184 588464 282236 588470
rect 282184 588406 282236 588412
rect 282920 588464 282972 588470
rect 282920 588406 282972 588412
rect 267004 579692 267056 579698
rect 267004 579634 267056 579640
rect 282196 575550 282224 588406
rect 280804 575544 280856 575550
rect 280804 575486 280856 575492
rect 282184 575544 282236 575550
rect 282184 575486 282236 575492
rect 280816 561746 280844 575486
rect 280804 561740 280856 561746
rect 280804 561682 280856 561688
rect 278044 561672 278096 561678
rect 278044 561614 278096 561620
rect 278056 523734 278084 561614
rect 414676 558890 414704 595070
rect 525076 562358 525104 614178
rect 525168 607170 525196 616762
rect 525156 607164 525208 607170
rect 525156 607106 525208 607112
rect 527640 607164 527692 607170
rect 527640 607106 527692 607112
rect 527652 603770 527680 607106
rect 527640 603764 527692 603770
rect 527640 603706 527692 603712
rect 533344 603764 533396 603770
rect 533344 603706 533396 603712
rect 533356 592006 533384 603706
rect 533344 592000 533396 592006
rect 533344 591942 533396 591948
rect 525064 562352 525116 562358
rect 525064 562294 525116 562300
rect 533344 562352 533396 562358
rect 533344 562294 533396 562300
rect 414664 558884 414716 558890
rect 414664 558826 414716 558832
rect 416044 558884 416096 558890
rect 416044 558826 416096 558832
rect 416056 529922 416084 558826
rect 533356 543862 533384 562294
rect 533344 543856 533396 543862
rect 533344 543798 533396 543804
rect 535736 543856 535788 543862
rect 535736 543798 535788 543804
rect 535748 542366 535776 543798
rect 535736 542360 535788 542366
rect 535736 542302 535788 542308
rect 538036 542360 538088 542366
rect 538036 542302 538088 542308
rect 416044 529916 416096 529922
rect 416044 529858 416096 529864
rect 417516 529916 417568 529922
rect 417516 529858 417568 529864
rect 417528 526318 417556 529858
rect 417516 526312 417568 526318
rect 417516 526254 417568 526260
rect 418896 526312 418948 526318
rect 418896 526254 418948 526260
rect 278044 523728 278096 523734
rect 278044 523670 278096 523676
rect 418908 521626 418936 526254
rect 418896 521620 418948 521626
rect 418896 521562 418948 521568
rect 420184 521620 420236 521626
rect 420184 521562 420236 521568
rect 420196 514758 420224 521562
rect 420184 514752 420236 514758
rect 420184 514694 420236 514700
rect 422944 514752 422996 514758
rect 422944 514694 422996 514700
rect 422956 505782 422984 514694
rect 422944 505776 422996 505782
rect 422944 505718 422996 505724
rect 424324 505776 424376 505782
rect 424324 505718 424376 505724
rect 424336 480962 424364 505718
rect 266360 480956 266412 480962
rect 266360 480898 266412 480904
rect 424324 480956 424376 480962
rect 424324 480898 424376 480904
rect 437388 480956 437440 480962
rect 437388 480898 437440 480904
rect 437400 479602 437428 480898
rect 240784 479596 240836 479602
rect 240784 479538 240836 479544
rect 437388 479596 437440 479602
rect 437388 479538 437440 479544
rect 240324 478916 240376 478922
rect 240324 478858 240376 478864
rect 300216 180260 300268 180266
rect 300216 180202 300268 180208
rect 373736 180254 373888 180282
rect 300124 180192 300176 180198
rect 300124 180134 300176 180140
rect 239864 178832 239916 178838
rect 239864 178774 239916 178780
rect 239680 178492 239732 178498
rect 239680 178434 239732 178440
rect 241992 177750 242020 180132
rect 241980 177744 242032 177750
rect 241980 177686 242032 177692
rect 245948 177342 245976 180132
rect 245936 177336 245988 177342
rect 245936 177278 245988 177284
rect 239036 177268 239088 177274
rect 239036 177210 239088 177216
rect 235264 175228 235316 175234
rect 235264 175170 235316 175176
rect 249904 161474 249932 180132
rect 249812 161446 249932 161474
rect 249812 60722 249840 161446
rect 249800 60716 249852 60722
rect 249800 60658 249852 60664
rect 253952 6798 253980 180132
rect 257908 174146 257936 180132
rect 256700 174140 256752 174146
rect 256700 174082 256752 174088
rect 257896 174140 257948 174146
rect 257896 174082 257948 174088
rect 256712 100706 256740 174082
rect 261956 161474 261984 180132
rect 265912 161474 265940 180132
rect 269960 161474 269988 180132
rect 273916 177206 273944 180132
rect 273904 177200 273956 177206
rect 273904 177142 273956 177148
rect 277964 161474 277992 180132
rect 280068 178832 280120 178838
rect 280068 178774 280120 178780
rect 280080 176254 280108 178774
rect 281920 177750 281948 180132
rect 282920 178764 282972 178770
rect 282920 178706 282972 178712
rect 281908 177744 281960 177750
rect 281908 177686 281960 177692
rect 282932 176322 282960 178706
rect 282920 176316 282972 176322
rect 282920 176258 282972 176264
rect 280068 176248 280120 176254
rect 280068 176190 280120 176196
rect 285968 161474 285996 180132
rect 289924 177954 289952 180132
rect 289912 177948 289964 177954
rect 289912 177890 289964 177896
rect 293972 177614 294000 180132
rect 297928 179926 297956 180132
rect 297916 179920 297968 179926
rect 297916 179862 297968 179868
rect 300136 177954 300164 180134
rect 300124 177948 300176 177954
rect 300124 177890 300176 177896
rect 300228 177750 300256 180202
rect 301990 180118 302280 180146
rect 305946 180118 306236 180146
rect 309994 180118 310376 180146
rect 313950 180118 314240 180146
rect 317998 180118 318288 180146
rect 321954 180118 322336 180146
rect 326002 180118 326384 180146
rect 329958 180118 330248 180146
rect 334006 180118 334296 180146
rect 337962 180118 338068 180146
rect 342010 180118 342208 180146
rect 345966 180118 346256 180146
rect 349922 180118 350304 180146
rect 353970 180118 354352 180146
rect 357926 180118 358216 180146
rect 361974 180118 362264 180146
rect 365930 180118 366312 180146
rect 369978 180118 370360 180146
rect 302252 179518 302280 180118
rect 302240 179512 302292 179518
rect 302240 179454 302292 179460
rect 300216 177744 300268 177750
rect 300216 177686 300268 177692
rect 306208 177682 306236 180118
rect 310348 179586 310376 180118
rect 310336 179580 310388 179586
rect 310336 179522 310388 179528
rect 310428 178764 310480 178770
rect 310428 178706 310480 178712
rect 306196 177676 306248 177682
rect 306196 177618 306248 177624
rect 310440 177614 310468 178706
rect 293960 177608 294012 177614
rect 293960 177550 294012 177556
rect 310428 177608 310480 177614
rect 310428 177550 310480 177556
rect 314212 177546 314240 180118
rect 318260 179654 318288 180118
rect 318248 179648 318300 179654
rect 318248 179590 318300 179596
rect 314200 177540 314252 177546
rect 314200 177482 314252 177488
rect 322308 177138 322336 180118
rect 322296 177132 322348 177138
rect 322296 177074 322348 177080
rect 326356 176458 326384 180118
rect 330220 176526 330248 180118
rect 334268 178022 334296 180118
rect 338040 179450 338068 180118
rect 338028 179444 338080 179450
rect 338028 179386 338080 179392
rect 334256 178016 334308 178022
rect 334256 177958 334308 177964
rect 342180 177750 342208 180118
rect 346228 179489 346256 180118
rect 346214 179480 346270 179489
rect 346214 179415 346270 179424
rect 342168 177744 342220 177750
rect 342168 177686 342220 177692
rect 350276 177614 350304 180118
rect 350264 177608 350316 177614
rect 350264 177550 350316 177556
rect 354324 177449 354352 180118
rect 355692 178832 355744 178838
rect 355692 178774 355744 178780
rect 355704 178022 355732 178774
rect 355692 178016 355744 178022
rect 355692 177958 355744 177964
rect 358188 177478 358216 180118
rect 358176 177472 358228 177478
rect 354310 177440 354366 177449
rect 358176 177414 358228 177420
rect 362236 177410 362264 180118
rect 366284 178566 366312 180118
rect 370332 179761 370360 180118
rect 370318 179752 370374 179761
rect 370318 179687 370374 179696
rect 373736 179081 373764 180254
rect 377982 180118 378088 180146
rect 381938 180118 382228 180146
rect 373722 179072 373778 179081
rect 373722 179007 373778 179016
rect 366272 178560 366324 178566
rect 366272 178502 366324 178508
rect 354310 177375 354366 177384
rect 362224 177404 362276 177410
rect 362224 177346 362276 177352
rect 330208 176520 330260 176526
rect 330208 176462 330260 176468
rect 326344 176452 326396 176458
rect 326344 176394 326396 176400
rect 378060 176390 378088 180118
rect 382200 177342 382228 180118
rect 385604 180118 385940 180146
rect 389942 180118 390232 180146
rect 382188 177336 382240 177342
rect 382188 177278 382240 177284
rect 378048 176384 378100 176390
rect 378048 176326 378100 176332
rect 385604 176322 385632 180118
rect 390204 179722 390232 180118
rect 393608 180118 393944 180146
rect 397946 180118 398328 180146
rect 390192 179716 390244 179722
rect 390192 179658 390244 179664
rect 393608 178498 393636 180118
rect 393596 178492 393648 178498
rect 393596 178434 393648 178440
rect 398300 176322 398328 180118
rect 401704 180118 401948 180146
rect 405752 180118 405904 180146
rect 409998 180118 410104 180146
rect 401600 178696 401652 178702
rect 401600 178638 401652 178644
rect 401612 177585 401640 178638
rect 401414 177576 401470 177585
rect 401414 177511 401470 177520
rect 401598 177576 401654 177585
rect 401598 177511 401654 177520
rect 401428 177426 401456 177511
rect 401704 177426 401732 180118
rect 401428 177398 401732 177426
rect 385592 176316 385644 176322
rect 385592 176258 385644 176264
rect 398288 176316 398340 176322
rect 398288 176258 398340 176264
rect 405752 176254 405780 180118
rect 408500 178696 408552 178702
rect 408500 178638 408552 178644
rect 406200 178084 406252 178090
rect 406200 178026 406252 178032
rect 406212 177206 406240 178026
rect 406200 177200 406252 177206
rect 406200 177142 406252 177148
rect 408512 177138 408540 178638
rect 410076 178634 410104 180118
rect 413572 180118 413908 180146
rect 417620 180118 417956 180146
rect 421576 180118 421912 180146
rect 425624 180118 425960 180146
rect 429580 180118 429916 180146
rect 433628 180118 433964 180146
rect 437584 180118 437920 180146
rect 441724 180118 441968 180146
rect 445772 180118 445924 180146
rect 449926 180118 450032 180146
rect 410064 178628 410116 178634
rect 410064 178570 410116 178576
rect 413572 177274 413600 180118
rect 413560 177268 413612 177274
rect 413560 177210 413612 177216
rect 408500 177132 408552 177138
rect 408500 177074 408552 177080
rect 417620 176497 417648 180118
rect 421576 177721 421604 180118
rect 421562 177712 421618 177721
rect 421562 177647 421618 177656
rect 425624 176594 425652 180118
rect 429580 179625 429608 180118
rect 429566 179616 429622 179625
rect 429566 179551 429622 179560
rect 433628 177857 433656 180118
rect 437584 178809 437612 180118
rect 437570 178800 437626 178809
rect 437570 178735 437626 178744
rect 433614 177848 433670 177857
rect 433614 177783 433670 177792
rect 441724 176633 441752 180118
rect 445772 178945 445800 180118
rect 450004 178974 450032 180118
rect 453592 180118 453928 180146
rect 457548 180118 457884 180146
rect 461596 180118 461932 180146
rect 465552 180118 465888 180146
rect 469600 180118 469936 180146
rect 473556 180118 473892 180146
rect 477604 180118 477940 180146
rect 481652 180118 481896 180146
rect 485792 180118 485944 180146
rect 489946 180118 490052 180146
rect 453592 179217 453620 180118
rect 453578 179208 453634 179217
rect 453578 179143 453634 179152
rect 449992 178968 450044 178974
rect 445758 178936 445814 178945
rect 449992 178910 450044 178916
rect 445758 178871 445814 178880
rect 449898 178664 449954 178673
rect 449898 178599 449954 178608
rect 449912 177449 449940 178599
rect 449898 177440 449954 177449
rect 449898 177375 449954 177384
rect 441710 176624 441766 176633
rect 425612 176588 425664 176594
rect 441710 176559 441766 176568
rect 425612 176530 425664 176536
rect 417606 176488 417662 176497
rect 417606 176423 417662 176432
rect 405740 176248 405792 176254
rect 405740 176190 405792 176196
rect 457548 175234 457576 180118
rect 461596 176662 461624 180118
rect 465552 177993 465580 180118
rect 469600 179353 469628 180118
rect 469586 179344 469642 179353
rect 469586 179279 469642 179288
rect 465538 177984 465594 177993
rect 465538 177919 465594 177928
rect 473556 177585 473584 180118
rect 477604 178906 477632 180118
rect 477592 178900 477644 178906
rect 477592 178842 477644 178848
rect 481652 177818 481680 180118
rect 485792 179246 485820 180118
rect 485780 179240 485832 179246
rect 485780 179182 485832 179188
rect 490024 177886 490052 180118
rect 493612 180118 493948 180146
rect 497568 180118 497904 180146
rect 501616 180118 501952 180146
rect 505572 180118 505908 180146
rect 509620 180118 509956 180146
rect 513576 180118 513912 180146
rect 517624 180118 517960 180146
rect 521672 180118 521916 180146
rect 525812 180118 525964 180146
rect 529966 180118 530072 180146
rect 493612 179314 493640 180118
rect 493600 179308 493652 179314
rect 493600 179250 493652 179256
rect 490012 177880 490064 177886
rect 490012 177822 490064 177828
rect 481640 177812 481692 177818
rect 481640 177754 481692 177760
rect 490564 177812 490616 177818
rect 490564 177754 490616 177760
rect 473542 177576 473598 177585
rect 473542 177511 473598 177520
rect 461584 176656 461636 176662
rect 461584 176598 461636 176604
rect 457536 175228 457588 175234
rect 457536 175170 457588 175176
rect 260852 161446 261984 161474
rect 264992 161446 265940 161474
rect 269132 161446 269988 161474
rect 277412 161446 277992 161474
rect 285692 161446 285996 161474
rect 256700 100700 256752 100706
rect 256700 100642 256752 100648
rect 260852 33114 260880 161446
rect 264992 139398 265020 161446
rect 264980 139392 265032 139398
rect 264980 139334 265032 139340
rect 269132 73166 269160 161446
rect 277412 113150 277440 161446
rect 285692 153202 285720 161446
rect 285680 153196 285732 153202
rect 285680 153138 285732 153144
rect 490576 150414 490604 177754
rect 497568 177002 497596 180118
rect 501616 179042 501644 180118
rect 501604 179036 501656 179042
rect 501604 178978 501656 178984
rect 505572 177070 505600 180118
rect 509620 179110 509648 180118
rect 509608 179104 509660 179110
rect 509608 179046 509660 179052
rect 513576 177818 513604 180118
rect 517624 179382 517652 180118
rect 517612 179376 517664 179382
rect 517612 179318 517664 179324
rect 521672 179178 521700 180118
rect 521660 179172 521712 179178
rect 521660 179114 521712 179120
rect 513564 177812 513616 177818
rect 513564 177754 513616 177760
rect 505560 177064 505612 177070
rect 505560 177006 505612 177012
rect 497556 176996 497608 177002
rect 497556 176938 497608 176944
rect 490564 150408 490616 150414
rect 490564 150350 490616 150356
rect 525812 137970 525840 180118
rect 530044 161474 530072 180118
rect 532712 180118 533968 180146
rect 536852 180118 537970 180146
rect 531964 178016 532016 178022
rect 531964 177958 532016 177964
rect 530676 177812 530728 177818
rect 530676 177754 530728 177760
rect 530688 176322 530716 177754
rect 531976 176390 532004 177958
rect 531964 176384 532016 176390
rect 531964 176326 532016 176332
rect 530676 176316 530728 176322
rect 530676 176258 530728 176264
rect 529952 161446 530072 161474
rect 525800 137964 525852 137970
rect 525800 137906 525852 137912
rect 277400 113144 277452 113150
rect 277400 113086 277452 113092
rect 529952 85542 529980 161446
rect 529940 85536 529992 85542
rect 529940 85478 529992 85484
rect 269120 73160 269172 73166
rect 269120 73102 269172 73108
rect 532712 45558 532740 180118
rect 532700 45552 532752 45558
rect 532700 45494 532752 45500
rect 260840 33108 260892 33114
rect 260840 33050 260892 33056
rect 536852 6866 536880 180118
rect 536932 179104 536984 179110
rect 536932 179046 536984 179052
rect 536944 177818 536972 179046
rect 538048 178022 538076 542302
rect 538036 178016 538088 178022
rect 538036 177958 538088 177964
rect 536932 177812 536984 177818
rect 536932 177754 536984 177760
rect 538232 177342 538260 700266
rect 538312 592000 538364 592006
rect 538312 591942 538364 591948
rect 538324 179722 538352 591942
rect 538404 479528 538456 479534
rect 538404 479470 538456 479476
rect 538312 179716 538364 179722
rect 538312 179658 538364 179664
rect 538416 179110 538444 479470
rect 538956 418192 539008 418198
rect 538956 418134 539008 418140
rect 538968 412634 538996 418134
rect 538876 412606 538996 412634
rect 538404 179104 538456 179110
rect 538404 179046 538456 179052
rect 538876 177546 538904 412606
rect 538956 364404 539008 364410
rect 538956 364346 539008 364352
rect 538968 177682 538996 364346
rect 540244 324352 540296 324358
rect 540244 324294 540296 324300
rect 540256 179654 540284 324294
rect 540336 271924 540388 271930
rect 540336 271866 540388 271872
rect 540244 179648 540296 179654
rect 540244 179590 540296 179596
rect 540348 179586 540376 271866
rect 540428 231872 540480 231878
rect 540428 231814 540480 231820
rect 540336 179580 540388 179586
rect 540336 179522 540388 179528
rect 540440 179518 540468 231814
rect 540428 179512 540480 179518
rect 540428 179454 540480 179460
rect 538956 177676 539008 177682
rect 538956 177618 539008 177624
rect 538864 177540 538916 177546
rect 538864 177482 538916 177488
rect 542372 177410 542400 702406
rect 580262 644056 580318 644065
rect 580262 643991 580318 644000
rect 579618 577688 579674 577697
rect 579618 577623 579674 577632
rect 579632 577250 579660 577623
rect 577504 577244 577556 577250
rect 577504 577186 577556 577192
rect 579620 577244 579672 577250
rect 579620 577186 579672 577192
rect 543004 378208 543056 378214
rect 543004 378150 543056 378156
rect 542360 177404 542412 177410
rect 542360 177346 542412 177352
rect 538220 177336 538272 177342
rect 538220 177278 538272 177284
rect 543016 176458 543044 378150
rect 577516 179450 577544 577186
rect 579618 524512 579674 524521
rect 577596 524476 577648 524482
rect 579618 524447 579620 524456
rect 577596 524418 577648 524424
rect 579672 524447 579674 524456
rect 579620 524418 579672 524424
rect 577504 179444 577556 179450
rect 577504 179386 577556 179392
rect 577608 176526 577636 524418
rect 579618 418296 579674 418305
rect 579618 418231 579674 418240
rect 579632 418198 579660 418231
rect 579620 418192 579672 418198
rect 579620 418134 579672 418140
rect 580170 378448 580226 378457
rect 580170 378383 580226 378392
rect 580184 378214 580212 378383
rect 580172 378208 580224 378214
rect 580172 378150 580224 378156
rect 580170 365120 580226 365129
rect 580170 365055 580226 365064
rect 580184 364410 580212 365055
rect 580172 364404 580224 364410
rect 580172 364346 580224 364352
rect 579618 325272 579674 325281
rect 579618 325207 579674 325216
rect 579632 324358 579660 325207
rect 579620 324352 579672 324358
rect 579620 324294 579672 324300
rect 580170 272232 580226 272241
rect 580170 272167 580226 272176
rect 580184 271930 580212 272167
rect 580172 271924 580224 271930
rect 580172 271866 580224 271872
rect 580170 232384 580226 232393
rect 580170 232319 580226 232328
rect 580184 231878 580212 232319
rect 580172 231872 580224 231878
rect 580172 231814 580224 231820
rect 580170 219056 580226 219065
rect 580170 218991 580226 219000
rect 580078 192536 580134 192545
rect 580078 192471 580134 192480
rect 580092 178770 580120 192471
rect 580184 180266 580212 218991
rect 580172 180260 580224 180266
rect 580172 180202 580224 180208
rect 580170 179208 580226 179217
rect 580170 179143 580226 179152
rect 580080 178764 580132 178770
rect 580080 178706 580132 178712
rect 580184 178090 580212 179143
rect 580276 178566 580304 643991
rect 580354 591016 580410 591025
rect 580354 590951 580410 590960
rect 580264 178560 580316 178566
rect 580264 178502 580316 178508
rect 580172 178084 580224 178090
rect 580172 178026 580224 178032
rect 580368 177478 580396 590951
rect 580446 537840 580502 537849
rect 580446 537775 580502 537784
rect 580460 177614 580488 537775
rect 580538 484664 580594 484673
rect 580538 484599 580594 484608
rect 580552 177750 580580 484599
rect 580630 471472 580686 471481
rect 580630 471407 580686 471416
rect 580644 178702 580672 471407
rect 580722 431624 580778 431633
rect 580722 431559 580778 431568
rect 580736 178838 580764 431559
rect 580814 312080 580870 312089
rect 580814 312015 580870 312024
rect 580828 180130 580856 312015
rect 580906 258904 580962 258913
rect 580906 258839 580962 258848
rect 580920 180198 580948 258839
rect 580908 180192 580960 180198
rect 580908 180134 580960 180140
rect 580816 180124 580868 180130
rect 580816 180066 580868 180072
rect 580724 178832 580776 178838
rect 580724 178774 580776 178780
rect 580632 178696 580684 178702
rect 580632 178638 580684 178644
rect 580540 177744 580592 177750
rect 580540 177686 580592 177692
rect 580448 177608 580500 177614
rect 580448 177550 580500 177556
rect 580356 177472 580408 177478
rect 580356 177414 580408 177420
rect 577596 176520 577648 176526
rect 577596 176462 577648 176468
rect 543004 176452 543056 176458
rect 543004 176394 543056 176400
rect 580172 153196 580224 153202
rect 580172 153138 580224 153144
rect 580184 152697 580212 153138
rect 580170 152688 580226 152697
rect 580170 152623 580226 152632
rect 580172 139392 580224 139398
rect 580170 139360 580172 139369
rect 580224 139360 580226 139369
rect 580170 139295 580226 139304
rect 579804 113144 579856 113150
rect 579804 113086 579856 113092
rect 579816 112849 579844 113086
rect 579802 112840 579858 112849
rect 579802 112775 579858 112784
rect 580172 100700 580224 100706
rect 580172 100642 580224 100648
rect 580184 99521 580212 100642
rect 580170 99512 580226 99521
rect 580170 99447 580226 99456
rect 580172 73160 580224 73166
rect 580172 73102 580224 73108
rect 580184 73001 580212 73102
rect 580170 72992 580226 73001
rect 580170 72927 580226 72936
rect 580172 60716 580224 60722
rect 580172 60658 580224 60664
rect 580184 59673 580212 60658
rect 580170 59664 580226 59673
rect 580170 59599 580226 59608
rect 580170 33144 580226 33153
rect 580170 33079 580172 33088
rect 580224 33079 580226 33088
rect 580172 33050 580224 33056
rect 536840 6860 536892 6866
rect 536840 6802 536892 6808
rect 253940 6792 253992 6798
rect 253940 6734 253992 6740
rect 580172 6792 580224 6798
rect 580172 6734 580224 6740
rect 580184 6633 580212 6734
rect 580170 6624 580226 6633
rect 580170 6559 580226 6568
rect 47584 3460 47636 3466
rect 47584 3402 47636 3408
rect 1646 354 1758 480
rect 1412 326 1758 354
rect 1646 -960 1758 326
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 8114 700304 8170 700360
rect 3422 671200 3478 671256
rect 3054 566888 3110 566944
rect 3330 514820 3386 514856
rect 3330 514800 3332 514820
rect 3332 514800 3384 514820
rect 3384 514800 3386 514820
rect 3330 501744 3386 501800
rect 3330 449520 3386 449576
rect 3330 397468 3332 397488
rect 3332 397468 3384 397488
rect 3384 397468 3386 397488
rect 3330 397432 3386 397468
rect 3054 345344 3110 345400
rect 3146 293120 3202 293176
rect 3238 241032 3294 241088
rect 3330 188808 3386 188864
rect 3514 658144 3570 658200
rect 3514 606056 3570 606112
rect 3422 177792 3478 177848
rect 3606 553832 3662 553888
rect 3606 462576 3662 462632
rect 3698 410488 3754 410544
rect 3790 358400 3846 358456
rect 3606 177928 3662 177984
rect 3882 306176 3938 306232
rect 3974 254088 4030 254144
rect 4066 201864 4122 201920
rect 137834 700576 137890 700632
rect 89166 700440 89222 700496
rect 151358 466248 151414 466304
rect 91190 465160 91246 465216
rect 93674 465180 93730 465216
rect 93674 465160 93676 465180
rect 93676 465160 93728 465180
rect 93728 465160 93730 465180
rect 157246 466384 157302 466440
rect 96158 465196 96160 465216
rect 96160 465196 96212 465216
rect 96212 465196 96214 465216
rect 96158 465160 96214 465196
rect 101310 465160 101366 465216
rect 103702 465160 103758 465216
rect 106186 465160 106242 465216
rect 108486 465160 108542 465216
rect 111062 465160 111118 465216
rect 128726 465160 128782 465216
rect 136086 465160 136142 465216
rect 141054 465160 141110 465216
rect 146022 465160 146078 465216
rect 154486 465160 154542 465216
rect 168470 465160 168526 465216
rect 169758 465160 169814 465216
rect 131118 463936 131174 463992
rect 83462 463664 83518 463720
rect 88522 463664 88578 463720
rect 98550 463664 98606 463720
rect 113638 463664 113694 463720
rect 116122 463664 116178 463720
rect 118606 463664 118662 463720
rect 120998 463664 121054 463720
rect 123574 463664 123630 463720
rect 125966 463664 126022 463720
rect 133510 463664 133566 463720
rect 138478 463664 138534 463720
rect 143630 463664 143686 463720
rect 148506 463664 148562 463720
rect 48042 416880 48098 416936
rect 47950 415928 48006 415984
rect 47582 388320 47638 388376
rect 47858 388048 47914 388104
rect 48226 413752 48282 413808
rect 48134 389952 48190 390008
rect 49330 412800 49386 412856
rect 49238 409944 49294 410000
rect 49422 411018 49478 411074
rect 49606 408162 49662 408218
rect 110970 379616 111026 379672
rect 113546 379616 113602 379672
rect 118330 379616 118386 379672
rect 120998 379616 121054 379672
rect 123482 379616 123538 379672
rect 130934 379616 130990 379672
rect 144918 379616 144974 379672
rect 87050 379480 87106 379536
rect 88154 379480 88210 379536
rect 89442 379480 89498 379536
rect 90730 379480 90786 379536
rect 116030 379500 116086 379536
rect 116030 379480 116032 379500
rect 116032 379480 116084 379500
rect 116084 379480 116086 379500
rect 150990 379480 151046 379536
rect 67546 377984 67602 378040
rect 74354 377984 74410 378040
rect 78494 377984 78550 378040
rect 81162 377984 81218 378040
rect 85946 377984 86002 378040
rect 91926 378020 91928 378040
rect 91928 378020 91980 378040
rect 91980 378020 91982 378040
rect 91926 377984 91982 378020
rect 92846 378004 92902 378040
rect 92846 377984 92848 378004
rect 92848 377984 92900 378004
rect 92900 377984 92902 378004
rect 66166 377032 66222 377088
rect 68926 377032 68982 377088
rect 70306 377032 70362 377088
rect 71686 377032 71742 377088
rect 73066 377032 73122 377088
rect 75826 377032 75882 377088
rect 77206 377032 77262 377088
rect 78310 377052 78366 377088
rect 78310 377032 78312 377052
rect 78312 377032 78364 377052
rect 78364 377032 78366 377052
rect 74446 376896 74502 376952
rect 79966 377032 80022 377088
rect 81254 377032 81310 377088
rect 82726 377032 82782 377088
rect 84106 377032 84162 377088
rect 85486 377032 85542 377088
rect 81346 376896 81402 376952
rect 84014 376896 84070 376952
rect 93950 377984 94006 378040
rect 95238 377984 95294 378040
rect 96526 377984 96582 378040
rect 97630 377984 97686 378040
rect 99930 377984 99986 378040
rect 104806 377984 104862 378040
rect 106094 377984 106150 378040
rect 108486 377984 108542 378040
rect 125966 377984 126022 378040
rect 128542 377984 128598 378040
rect 133510 377984 133566 378040
rect 96434 377848 96490 377904
rect 86774 377032 86830 377088
rect 89626 377032 89682 377088
rect 92386 377032 92442 377088
rect 93766 377032 93822 377088
rect 102046 377712 102102 377768
rect 99286 377032 99342 377088
rect 140778 378664 140834 378720
rect 136086 377984 136142 378040
rect 138662 377984 138718 378040
rect 141146 377984 141202 378040
rect 146022 377984 146078 378040
rect 148598 377984 148654 378040
rect 153382 377984 153438 378040
rect 155958 377984 156014 378040
rect 180706 377304 180762 377360
rect 173806 377168 173862 377224
rect 173714 376896 173770 376952
rect 117226 286492 117228 286512
rect 117228 286492 117280 286512
rect 117280 286492 117282 286512
rect 117226 286456 117282 286492
rect 48134 236816 48190 236872
rect 47950 235864 48006 235920
rect 47766 232736 47822 232792
rect 47674 230968 47730 231024
rect 47858 229880 47914 229936
rect 47766 199688 47822 199744
rect 47674 199552 47730 199608
rect 48042 233688 48098 233744
rect 47858 197240 47914 197296
rect 49514 228162 49570 228218
rect 49330 209888 49386 209944
rect 48134 199824 48190 199880
rect 49422 208034 49478 208090
rect 108946 285948 108948 285968
rect 108948 285948 109000 285968
rect 109000 285948 109002 285968
rect 108946 285912 109002 285948
rect 111706 285912 111762 285968
rect 136546 286356 136548 286376
rect 136548 286356 136600 286376
rect 136600 286356 136602 286376
rect 136546 286320 136602 286356
rect 126886 286084 126888 286104
rect 126888 286084 126940 286104
rect 126940 286084 126942 286104
rect 126886 286048 126942 286084
rect 132314 286048 132370 286104
rect 133786 286048 133842 286104
rect 79966 285676 79968 285696
rect 79968 285676 80020 285696
rect 80020 285676 80022 285696
rect 79966 285640 80022 285676
rect 81346 285640 81402 285696
rect 86866 285640 86922 285696
rect 89626 285640 89682 285696
rect 93674 285640 93730 285696
rect 102046 285640 102102 285696
rect 104806 285640 104862 285696
rect 106186 285640 106242 285696
rect 121366 285640 121422 285696
rect 96158 285096 96214 285152
rect 113822 285096 113878 285152
rect 123574 285132 123576 285152
rect 123576 285132 123628 285152
rect 123628 285132 123630 285152
rect 123574 285096 123630 285132
rect 128726 285096 128782 285152
rect 98550 284996 98552 285016
rect 98552 284996 98604 285016
rect 98604 284996 98606 285016
rect 98550 284960 98606 284996
rect 118606 284960 118662 285016
rect 91190 284824 91246 284880
rect 169666 286184 169722 286240
rect 139306 285640 139362 285696
rect 142066 285640 142122 285696
rect 144826 285640 144882 285696
rect 146206 285640 146262 285696
rect 148966 285640 149022 285696
rect 151726 285640 151782 285696
rect 154486 285640 154542 285696
rect 157246 285640 157302 285696
rect 170678 286320 170734 286376
rect 189078 459176 189134 459232
rect 189078 399336 189134 399392
rect 189078 397704 189134 397760
rect 189078 396344 189134 396400
rect 189446 394848 189502 394904
rect 189078 393624 189134 393680
rect 180706 284008 180762 284064
rect 49606 208306 49662 208362
rect 70582 199416 70638 199472
rect 77758 199416 77814 199472
rect 78862 199416 78918 199472
rect 88614 199416 88670 199472
rect 91190 199416 91246 199472
rect 103702 199416 103758 199472
rect 111062 199416 111118 199472
rect 71870 198600 71926 198656
rect 75550 198600 75606 198656
rect 76838 198600 76894 198656
rect 80150 198600 80206 198656
rect 81346 198600 81402 198656
rect 82542 198600 82598 198656
rect 84566 198600 84622 198656
rect 86222 198636 86224 198656
rect 86224 198636 86276 198656
rect 86276 198636 86278 198656
rect 86222 198600 86278 198636
rect 87970 198600 88026 198656
rect 92846 198600 92902 198656
rect 93582 198600 93638 198656
rect 95974 198600 96030 198656
rect 104438 198600 104494 198656
rect 105910 198620 105966 198656
rect 105910 198600 105912 198620
rect 105912 198600 105964 198620
rect 105964 198600 105966 198620
rect 73434 198328 73490 198384
rect 67546 198192 67602 198248
rect 66166 197376 66222 197432
rect 69662 197920 69718 197976
rect 68926 197376 68982 197432
rect 74354 198192 74410 198248
rect 83646 198192 83702 198248
rect 78586 197376 78642 197432
rect 81254 197376 81310 197432
rect 85854 198464 85910 198520
rect 88246 198464 88302 198520
rect 89534 198464 89590 198520
rect 90822 198464 90878 198520
rect 98366 198464 98422 198520
rect 100022 198464 100078 198520
rect 100942 198464 100998 198520
rect 102230 198464 102286 198520
rect 103334 198464 103390 198520
rect 100022 196832 100078 196888
rect 103334 196968 103390 197024
rect 102230 196696 102286 196752
rect 106094 198600 106150 198656
rect 108486 198600 108542 198656
rect 113638 198600 113694 198656
rect 117042 198600 117098 198656
rect 118422 198600 118478 198656
rect 107014 197920 107070 197976
rect 108578 197920 108634 197976
rect 109222 197920 109278 197976
rect 104438 196560 104494 196616
rect 120998 198636 121000 198656
rect 121000 198636 121052 198656
rect 121052 198636 121054 198656
rect 120998 198600 121054 198636
rect 123574 198600 123630 198656
rect 126610 198600 126666 198656
rect 128910 198600 128966 198656
rect 146022 198600 146078 198656
rect 153382 198600 153438 198656
rect 173438 198600 173494 198656
rect 138662 197784 138718 197840
rect 141238 197784 141294 197840
rect 143446 197784 143502 197840
rect 133510 197648 133566 197704
rect 148598 197648 148654 197704
rect 150990 197648 151046 197704
rect 173254 197784 173310 197840
rect 155958 197376 156014 197432
rect 189078 279112 189134 279168
rect 189078 219272 189134 219328
rect 189078 217640 189134 217696
rect 189170 216280 189226 216336
rect 189078 213696 189134 213752
rect 189630 199552 189686 199608
rect 189078 197240 189134 197296
rect 3422 149776 3478 149832
rect 3238 136720 3294 136776
rect 3146 84632 3202 84688
rect 3422 45500 3424 45520
rect 3424 45500 3476 45520
rect 3476 45500 3478 45520
rect 3422 45464 3478 45500
rect 3422 6432 3478 6488
rect 189814 465432 189870 465488
rect 189998 378936 190054 378992
rect 189814 198872 189870 198928
rect 190458 214784 190514 214840
rect 190366 199688 190422 199744
rect 191194 199008 191250 199064
rect 201498 177656 201554 177712
rect 235170 377712 235226 377768
rect 232870 198736 232926 198792
rect 232778 196832 232834 196888
rect 234986 197104 235042 197160
rect 235170 196696 235226 196752
rect 218058 177520 218114 177576
rect 237378 478916 237434 478952
rect 237378 478896 237380 478916
rect 237380 478896 237432 478916
rect 237432 478896 237434 478916
rect 237378 477808 237434 477864
rect 235354 465568 235410 465624
rect 237378 476720 237434 476776
rect 237378 473728 237434 473784
rect 237470 472640 237526 472696
rect 237378 472096 237434 472152
rect 235630 379072 235686 379128
rect 237378 469260 237434 469296
rect 237378 469240 237380 469260
rect 237380 469240 237432 469260
rect 237432 469240 237434 469260
rect 237378 467900 237434 467936
rect 237378 467880 237380 467900
rect 237380 467880 237432 467900
rect 237432 467880 237434 467900
rect 237378 466656 237434 466712
rect 237378 464752 237434 464808
rect 237378 462576 237434 462632
rect 237470 459448 237526 459504
rect 237378 458244 237434 458280
rect 237378 458224 237380 458244
rect 237380 458224 237432 458244
rect 237432 458224 237434 458244
rect 237378 449520 237434 449576
rect 237378 447344 237434 447400
rect 237378 444216 237434 444272
rect 237378 442312 237434 442368
rect 237378 439456 237434 439512
rect 237378 437552 237434 437608
rect 238022 454688 238078 454744
rect 238022 452648 238078 452704
rect 237930 434288 237986 434344
rect 237378 432112 237434 432168
rect 237378 431160 237434 431216
rect 237470 427080 237526 427136
rect 237378 426672 237434 426728
rect 237378 423580 237380 423600
rect 237380 423580 237432 423600
rect 237432 423580 237434 423600
rect 237378 423544 237434 423580
rect 237378 422340 237434 422376
rect 237378 422320 237380 422340
rect 237380 422320 237432 422340
rect 237432 422320 237434 422340
rect 237378 419192 237434 419248
rect 237378 416880 237434 416936
rect 237378 415928 237434 415984
rect 237378 413924 237380 413944
rect 237380 413924 237432 413944
rect 237432 413924 237434 413944
rect 237378 413888 237434 413924
rect 237378 411848 237434 411904
rect 237930 411304 237986 411360
rect 237378 408468 237434 408504
rect 237378 408448 237380 408468
rect 237380 408448 237432 408468
rect 237432 408448 237434 408468
rect 237838 407088 237894 407144
rect 237378 405748 237434 405784
rect 237378 405728 237380 405748
rect 237380 405728 237432 405748
rect 237432 405728 237434 405748
rect 237378 401784 237434 401840
rect 237378 400696 237434 400752
rect 237470 396616 237526 396672
rect 237378 396208 237434 396264
rect 237378 392128 237434 392184
rect 237378 390632 237434 390688
rect 237378 388728 237434 388784
rect 237378 386552 237434 386608
rect 237378 385464 237434 385520
rect 237378 383596 237380 383616
rect 237380 383596 237432 383616
rect 237432 383596 237434 383616
rect 237378 383560 237434 383596
rect 237470 381520 237526 381576
rect 237378 380976 237434 381032
rect 238298 446392 238354 446448
rect 238206 398792 238262 398848
rect 238114 393896 238170 393952
rect 237378 378020 237380 378040
rect 237380 378020 237432 378040
rect 237432 378020 237434 378040
rect 237378 377984 237434 378020
rect 235814 377576 235870 377632
rect 237378 377168 237434 377224
rect 238482 441632 238538 441688
rect 238390 403960 238446 404016
rect 238574 436192 238630 436248
rect 238482 379344 238538 379400
rect 238666 429120 238722 429176
rect 238666 420960 238722 421016
rect 238666 378664 238722 378720
rect 238298 377032 238354 377088
rect 237378 376660 237380 376680
rect 237380 376660 237432 376680
rect 237432 376660 237434 376680
rect 237378 376624 237434 376660
rect 237378 373632 237434 373688
rect 237378 372408 237434 372464
rect 237378 371048 237434 371104
rect 237378 368328 237434 368384
rect 237378 366988 237434 367024
rect 237378 366968 237380 366988
rect 237380 366968 237432 366988
rect 237432 366968 237434 366988
rect 237470 366424 237526 366480
rect 237378 362788 237380 362808
rect 237380 362788 237432 362808
rect 237432 362788 237434 362808
rect 237378 362752 237434 362788
rect 237470 362480 237526 362536
rect 237378 361392 237434 361448
rect 237378 360032 237434 360088
rect 237378 358708 237380 358728
rect 237380 358708 237432 358728
rect 237432 358708 237434 358728
rect 237378 358672 237434 358708
rect 237470 358400 237526 358456
rect 237378 357348 237380 357368
rect 237380 357348 237432 357368
rect 237432 357348 237434 357368
rect 237378 357312 237434 357348
rect 237378 355816 237434 355872
rect 237470 355272 237526 355328
rect 237378 354320 237434 354376
rect 237378 352960 237434 353016
rect 237378 351772 237380 351792
rect 237380 351772 237432 351792
rect 237432 351772 237434 351792
rect 237378 351736 237434 351772
rect 237470 351328 237526 351384
rect 237378 350240 237434 350296
rect 237378 349052 237380 349072
rect 237380 349052 237432 349072
rect 237432 349052 237434 349072
rect 237378 349016 237434 349052
rect 237470 347676 237526 347712
rect 237470 347656 237472 347676
rect 237472 347656 237524 347676
rect 237524 347656 237526 347676
rect 237378 347248 237434 347304
rect 237378 346160 237434 346216
rect 237378 344800 237434 344856
rect 238022 343576 238078 343632
rect 237378 343168 237434 343224
rect 237378 342080 237434 342136
rect 237378 340720 237434 340776
rect 237470 340176 237526 340232
rect 238114 339088 238170 339144
rect 237378 338036 237380 338056
rect 237380 338036 237432 338056
rect 237432 338036 237434 338056
rect 237378 338000 237434 338036
rect 237378 336504 237434 336560
rect 237470 336096 237526 336152
rect 237378 335008 237434 335064
rect 237378 333784 237434 333840
rect 237378 332424 237434 332480
rect 237470 332016 237526 332072
rect 237378 331064 237434 331120
rect 237378 329568 237434 329624
rect 237470 329024 237526 329080
rect 237378 327936 237434 327992
rect 237378 327020 237380 327040
rect 237380 327020 237432 327040
rect 237432 327020 237434 327040
rect 237378 326984 237434 327020
rect 237378 325488 237434 325544
rect 237378 324944 237434 325000
rect 237378 323856 237434 323912
rect 237470 322768 237526 322824
rect 237378 321444 237380 321464
rect 237380 321444 237432 321464
rect 237432 321444 237434 321464
rect 237378 321408 237434 321444
rect 237470 320864 237526 320920
rect 237378 319912 237434 319968
rect 237378 317364 237380 317384
rect 237380 317364 237432 317384
rect 237432 317364 237434 317384
rect 237378 317328 237434 317364
rect 237562 316784 237618 316840
rect 237378 315832 237434 315888
rect 237378 314472 237434 314528
rect 237378 313112 237434 313168
rect 237470 312704 237526 312760
rect 237378 311788 237380 311808
rect 237380 311788 237432 311808
rect 237432 311788 237434 311808
rect 237378 311752 237434 311788
rect 237378 309440 237434 309496
rect 237470 309204 237472 309224
rect 237472 309204 237524 309224
rect 237524 309204 237526 309224
rect 237470 309168 237526 309204
rect 237378 307828 237434 307864
rect 237378 307808 237380 307828
rect 237380 307808 237432 307828
rect 237432 307808 237434 307828
rect 238022 306448 238078 306504
rect 237470 305496 237526 305552
rect 237378 304988 237380 305008
rect 237380 304988 237432 305008
rect 237432 304988 237434 305008
rect 237378 304952 237434 304988
rect 237378 303864 237434 303920
rect 237378 302368 237434 302424
rect 237470 301416 237526 301472
rect 237378 300892 237434 300928
rect 237378 300872 237380 300892
rect 237380 300872 237432 300892
rect 237432 300872 237434 300892
rect 236734 300056 236790 300112
rect 235814 199824 235870 199880
rect 235906 196968 235962 197024
rect 235722 196560 235778 196616
rect 237378 298832 237434 298888
rect 237378 297880 237434 297936
rect 236826 296928 236882 296984
rect 237378 295840 237434 295896
rect 237378 294888 237434 294944
rect 236918 293800 236974 293856
rect 237378 292848 237434 292904
rect 237378 291760 237434 291816
rect 237010 290808 237066 290864
rect 237378 289876 237434 289912
rect 237378 289856 237380 289876
rect 237380 289856 237432 289876
rect 237432 289856 237434 289876
rect 237378 288768 237434 288824
rect 237102 287680 237158 287736
rect 237470 286728 237526 286784
rect 237378 285912 237434 285968
rect 237378 284688 237434 284744
rect 237470 283736 237526 283792
rect 237378 282820 237380 282840
rect 237380 282820 237432 282840
rect 237432 282820 237434 282840
rect 237378 282784 237434 282820
rect 237378 281696 237434 281752
rect 237470 280608 237526 280664
rect 237378 279792 237434 279848
rect 237470 275576 237526 275632
rect 237378 274780 237434 274816
rect 237378 274760 237380 274780
rect 237380 274760 237432 274780
rect 237432 274760 237434 274780
rect 237378 273672 237434 273728
rect 237378 272584 237434 272640
rect 237378 269456 237434 269512
rect 237378 265512 237434 265568
rect 237378 263472 237434 263528
rect 237470 260344 237526 260400
rect 237378 259548 237434 259584
rect 237378 259528 237380 259548
rect 237380 259528 237432 259548
rect 237432 259528 237434 259548
rect 237378 258440 237434 258496
rect 237378 256264 237434 256320
rect 237470 255448 237526 255504
rect 237378 254360 237434 254416
rect 237470 253272 237526 253328
rect 237378 252492 237380 252512
rect 237380 252492 237432 252512
rect 237432 252492 237434 252512
rect 237378 252456 237434 252492
rect 237378 250280 237434 250336
rect 237378 247288 237434 247344
rect 237378 246200 237434 246256
rect 237378 245112 237434 245168
rect 237378 242256 237434 242312
rect 237378 240216 237434 240272
rect 237378 237224 237434 237280
rect 237378 236020 237434 236056
rect 237378 236000 237380 236020
rect 237380 236000 237432 236020
rect 237432 236000 237434 236020
rect 237378 230968 237434 231024
rect 237470 228928 237526 228984
rect 237378 227976 237434 228032
rect 237378 227024 237434 227080
rect 237378 225936 237434 225992
rect 237378 223896 237434 223952
rect 237930 222944 237986 223000
rect 237378 221992 237434 222048
rect 237378 220904 237434 220960
rect 237378 218864 237434 218920
rect 237378 217776 237434 217832
rect 237378 215736 237434 215792
rect 237470 214784 237526 214840
rect 237378 213868 237380 213888
rect 237380 213868 237432 213888
rect 237432 213868 237434 213888
rect 237378 213832 237434 213868
rect 237378 212744 237434 212800
rect 237470 211928 237526 211984
rect 237470 210704 237526 210760
rect 237378 209788 237380 209808
rect 237380 209788 237432 209808
rect 237432 209788 237434 209808
rect 237378 209752 237434 209788
rect 237470 208800 237526 208856
rect 237378 207712 237434 207768
rect 237378 206624 237434 206680
rect 237470 205808 237526 205864
rect 237838 203632 237894 203688
rect 237378 202680 237434 202736
rect 237378 201592 237434 201648
rect 237378 200640 237434 200696
rect 237470 198600 237526 198656
rect 237378 197648 237434 197704
rect 237378 196696 237434 196752
rect 238114 270680 238170 270736
rect 238114 266464 238170 266520
rect 238022 216960 238078 217016
rect 238022 204584 238078 204640
rect 238298 278568 238354 278624
rect 238206 261568 238262 261624
rect 238206 257352 238262 257408
rect 238390 264560 238446 264616
rect 238390 251232 238446 251288
rect 238298 222808 238354 222864
rect 238298 219816 238354 219872
rect 238666 276800 238722 276856
rect 238574 267552 238630 267608
rect 238574 241168 238630 241224
rect 238482 232192 238538 232248
rect 238482 230016 238538 230072
rect 238666 224984 238722 225040
rect 237378 195608 237434 195664
rect 237470 194656 237526 194712
rect 237378 193568 237434 193624
rect 237378 192616 237434 192672
rect 237378 191528 237434 191584
rect 237470 190576 237526 190632
rect 237378 189624 237434 189680
rect 238390 188536 238446 188592
rect 238390 187604 238446 187640
rect 238390 187584 238392 187604
rect 238392 187584 238444 187604
rect 238444 187584 238446 187604
rect 238758 186496 238814 186552
rect 238022 185544 238078 185600
rect 238758 184456 238814 184512
rect 238390 183404 238392 183424
rect 238392 183404 238444 183424
rect 238444 183404 238446 183424
rect 238390 183368 238446 183404
rect 238298 182416 238354 182472
rect 238574 180512 238630 180568
rect 239402 181464 239458 181520
rect 239586 179152 239642 179208
rect 239310 178744 239366 178800
rect 239770 179288 239826 179344
rect 522854 596808 522910 596864
rect 346214 179424 346270 179480
rect 354310 177384 354366 177440
rect 370318 179696 370374 179752
rect 373722 179016 373778 179072
rect 401414 177520 401470 177576
rect 401598 177520 401654 177576
rect 421562 177656 421618 177712
rect 429566 179560 429622 179616
rect 437570 178744 437626 178800
rect 433614 177792 433670 177848
rect 453578 179152 453634 179208
rect 445758 178880 445814 178936
rect 449898 178608 449954 178664
rect 449898 177384 449954 177440
rect 441710 176568 441766 176624
rect 417606 176432 417662 176488
rect 469586 179288 469642 179344
rect 465538 177928 465594 177984
rect 473542 177520 473598 177576
rect 580262 644000 580318 644056
rect 579618 577632 579674 577688
rect 579618 524476 579674 524512
rect 579618 524456 579620 524476
rect 579620 524456 579672 524476
rect 579672 524456 579674 524476
rect 579618 418240 579674 418296
rect 580170 378392 580226 378448
rect 580170 365064 580226 365120
rect 579618 325216 579674 325272
rect 580170 272176 580226 272232
rect 580170 232328 580226 232384
rect 580170 219000 580226 219056
rect 580078 192480 580134 192536
rect 580170 179152 580226 179208
rect 580354 590960 580410 591016
rect 580446 537784 580502 537840
rect 580538 484608 580594 484664
rect 580630 471416 580686 471472
rect 580722 431568 580778 431624
rect 580814 312024 580870 312080
rect 580906 258848 580962 258904
rect 580170 152632 580226 152688
rect 580170 139340 580172 139360
rect 580172 139340 580224 139360
rect 580224 139340 580226 139360
rect 580170 139304 580226 139340
rect 579802 112784 579858 112840
rect 580170 99456 580226 99512
rect 580170 72936 580226 72992
rect 580170 59608 580226 59664
rect 580170 33108 580226 33144
rect 580170 33088 580172 33108
rect 580172 33088 580224 33108
rect 580224 33088 580226 33108
rect 580170 6568 580226 6624
<< metal3 >>
rect 137829 700634 137895 700637
rect 237966 700634 237972 700636
rect 137829 700632 237972 700634
rect 137829 700576 137834 700632
rect 137890 700576 237972 700632
rect 137829 700574 237972 700576
rect 137829 700571 137895 700574
rect 237966 700572 237972 700574
rect 238036 700572 238042 700636
rect 89161 700498 89227 700501
rect 235206 700498 235212 700500
rect 89161 700496 235212 700498
rect 89161 700440 89166 700496
rect 89222 700440 235212 700496
rect 89161 700438 235212 700440
rect 89161 700435 89227 700438
rect 235206 700436 235212 700438
rect 235276 700436 235282 700500
rect 8109 700362 8175 700365
rect 239254 700362 239260 700364
rect 8109 700360 239260 700362
rect 8109 700304 8114 700360
rect 8170 700304 239260 700360
rect 8109 700302 239260 700304
rect 8109 700299 8175 700302
rect 239254 700300 239260 700302
rect 239324 700300 239330 700364
rect -960 697220 480 697460
rect 580206 697172 580212 697236
rect 580276 697234 580282 697236
rect 583520 697234 584960 697324
rect 580276 697174 584960 697234
rect 580276 697172 580282 697174
rect 583520 697084 584960 697174
rect -960 684164 480 684404
rect 580390 683844 580396 683908
rect 580460 683906 580466 683908
rect 583520 683906 584960 683996
rect 580460 683846 584960 683906
rect 580460 683844 580466 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3417 671258 3483 671261
rect -960 671256 3483 671258
rect -960 671200 3422 671256
rect 3478 671200 3483 671256
rect -960 671198 3483 671200
rect -960 671108 480 671198
rect 3417 671195 3483 671198
rect 583520 670564 584960 670804
rect -960 658202 480 658292
rect 3509 658202 3575 658205
rect -960 658200 3575 658202
rect -960 658144 3514 658200
rect 3570 658144 3575 658200
rect -960 658142 3575 658144
rect -960 658052 480 658142
rect 3509 658139 3575 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 580257 644058 580323 644061
rect 583520 644058 584960 644148
rect 580257 644056 584960 644058
rect 580257 644000 580262 644056
rect 580318 644000 584960 644056
rect 580257 643998 584960 644000
rect 580257 643995 580323 643998
rect 583520 643908 584960 643998
rect -960 631940 480 632180
rect 580574 630804 580580 630868
rect 580644 630866 580650 630868
rect 583520 630866 584960 630956
rect 580644 630806 584960 630866
rect 580644 630804 580650 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect -960 619110 674 619170
rect -960 619034 480 619110
rect 614 619034 674 619110
rect -960 619020 674 619034
rect 246 618974 674 619020
rect 246 618490 306 618974
rect 246 618430 6930 618490
rect 6870 618354 6930 618430
rect 235390 618354 235396 618356
rect 6870 618294 235396 618354
rect 235390 618292 235396 618294
rect 235460 618292 235466 618356
rect 583520 617388 584960 617628
rect -960 606114 480 606204
rect 3509 606114 3575 606117
rect -960 606112 3575 606114
rect -960 606056 3514 606112
rect 3570 606056 3575 606112
rect -960 606054 3575 606056
rect -960 605964 480 606054
rect 3509 606051 3575 606054
rect 583520 604060 584960 604300
rect 522849 596866 522915 596869
rect 536782 596866 536788 596868
rect 522849 596864 536788 596866
rect 522849 596808 522854 596864
rect 522910 596808 536788 596864
rect 522849 596806 536788 596808
rect 522849 596803 522915 596806
rect 536782 596804 536788 596806
rect 536852 596804 536858 596868
rect -960 592908 480 593148
rect 580349 591018 580415 591021
rect 583520 591018 584960 591108
rect 580349 591016 584960 591018
rect 580349 590960 580354 591016
rect 580410 590960 584960 591016
rect 580349 590958 584960 590960
rect 580349 590955 580415 590958
rect 583520 590868 584960 590958
rect -960 579852 480 580092
rect 579613 577690 579679 577693
rect 583520 577690 584960 577780
rect 579613 577688 584960 577690
rect 579613 577632 579618 577688
rect 579674 577632 584960 577688
rect 579613 577630 584960 577632
rect 579613 577627 579679 577630
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 3049 566946 3115 566949
rect -960 566944 3115 566946
rect -960 566888 3054 566944
rect 3110 566888 3115 566944
rect -960 566886 3115 566888
rect -960 566796 480 566886
rect 3049 566883 3115 566886
rect 583520 564212 584960 564452
rect -960 553890 480 553980
rect 3601 553890 3667 553893
rect -960 553888 3667 553890
rect -960 553832 3606 553888
rect 3662 553832 3667 553888
rect -960 553830 3667 553832
rect -960 553740 480 553830
rect 3601 553827 3667 553830
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 580441 537842 580507 537845
rect 583520 537842 584960 537932
rect 580441 537840 584960 537842
rect 580441 537784 580446 537840
rect 580502 537784 584960 537840
rect 580441 537782 584960 537784
rect 580441 537779 580507 537782
rect 583520 537692 584960 537782
rect -960 527764 480 528004
rect 579613 524514 579679 524517
rect 583520 524514 584960 524604
rect 579613 524512 584960 524514
rect 579613 524456 579618 524512
rect 579674 524456 584960 524512
rect 579613 524454 584960 524456
rect 579613 524451 579679 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 3325 514858 3391 514861
rect -960 514856 3391 514858
rect -960 514800 3330 514856
rect 3386 514800 3391 514856
rect -960 514798 3391 514800
rect -960 514708 480 514798
rect 3325 514795 3391 514798
rect 583520 511172 584960 511412
rect -960 501802 480 501892
rect 3325 501802 3391 501805
rect -960 501800 3391 501802
rect -960 501744 3330 501800
rect 3386 501744 3391 501800
rect -960 501742 3391 501744
rect -960 501652 480 501742
rect 3325 501739 3391 501742
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 580533 484666 580599 484669
rect 583520 484666 584960 484756
rect 580533 484664 584960 484666
rect 580533 484608 580538 484664
rect 580594 484608 584960 484664
rect 580533 484606 584960 484608
rect 580533 484603 580599 484606
rect 583520 484516 584960 484606
rect 237373 478954 237439 478957
rect 240182 478954 240242 479400
rect 237373 478952 240242 478954
rect 237373 478896 237378 478952
rect 237434 478896 240242 478952
rect 237373 478894 240242 478896
rect 237373 478891 237439 478894
rect 237373 477866 237439 477869
rect 240182 477866 240242 478448
rect 237373 477864 240242 477866
rect 237373 477808 237378 477864
rect 237434 477808 240242 477864
rect 237373 477806 240242 477808
rect 237373 477803 237439 477806
rect 237373 476778 237439 476781
rect 240182 476778 240242 477360
rect 237373 476776 240242 476778
rect 237373 476720 237378 476776
rect 237434 476720 240242 476776
rect 237373 476718 240242 476720
rect 237373 476715 237439 476718
rect -960 475540 480 475780
rect 237373 473786 237439 473789
rect 240182 473786 240242 474368
rect 237373 473784 240242 473786
rect 237373 473728 237378 473784
rect 237434 473728 240242 473784
rect 237373 473726 240242 473728
rect 237373 473723 237439 473726
rect 237465 472698 237531 472701
rect 240182 472698 240242 473280
rect 237465 472696 240242 472698
rect 237465 472640 237470 472696
rect 237526 472640 240242 472696
rect 237465 472638 240242 472640
rect 237465 472635 237531 472638
rect 237373 472154 237439 472157
rect 240182 472154 240242 472328
rect 237373 472152 240242 472154
rect 237373 472096 237378 472152
rect 237434 472096 240242 472152
rect 237373 472094 240242 472096
rect 237373 472091 237439 472094
rect 580625 471474 580691 471477
rect 583520 471474 584960 471564
rect 580625 471472 584960 471474
rect 580625 471416 580630 471472
rect 580686 471416 584960 471472
rect 580625 471414 584960 471416
rect 580625 471411 580691 471414
rect 583520 471324 584960 471414
rect 237373 469298 237439 469301
rect 240182 469298 240242 469336
rect 237373 469296 240242 469298
rect 237373 469240 237378 469296
rect 237434 469240 240242 469296
rect 237373 469238 240242 469240
rect 237373 469235 237439 469238
rect 237373 467938 237439 467941
rect 240182 467938 240242 468248
rect 237373 467936 240242 467938
rect 237373 467880 237378 467936
rect 237434 467880 240242 467936
rect 237373 467878 240242 467880
rect 237373 467875 237439 467878
rect 237373 466714 237439 466717
rect 240182 466714 240242 467296
rect 237373 466712 240242 466714
rect 237373 466656 237378 466712
rect 237434 466656 240242 466712
rect 237373 466654 240242 466656
rect 237373 466651 237439 466654
rect 156086 466380 156092 466444
rect 156156 466442 156162 466444
rect 157241 466442 157307 466445
rect 156156 466440 157307 466442
rect 156156 466384 157246 466440
rect 157302 466384 157307 466440
rect 156156 466382 157307 466384
rect 156156 466380 156162 466382
rect 157241 466379 157307 466382
rect 151118 466244 151124 466308
rect 151188 466306 151194 466308
rect 151353 466306 151419 466309
rect 151188 466304 151419 466306
rect 151188 466248 151358 466304
rect 151414 466248 151419 466304
rect 151188 466246 151419 466248
rect 151188 466244 151194 466246
rect 151353 466243 151419 466246
rect 81014 465564 81020 465628
rect 81084 465626 81090 465628
rect 235349 465626 235415 465629
rect 81084 465624 235415 465626
rect 81084 465568 235354 465624
rect 235410 465568 235415 465624
rect 81084 465566 235415 465568
rect 81084 465564 81090 465566
rect 235349 465563 235415 465566
rect 86166 465428 86172 465492
rect 86236 465490 86242 465492
rect 189809 465490 189875 465493
rect 86236 465488 189875 465490
rect 86236 465432 189814 465488
rect 189870 465432 189875 465488
rect 86236 465430 189875 465432
rect 86236 465428 86242 465430
rect 189809 465427 189875 465430
rect 78806 465292 78812 465356
rect 78876 465354 78882 465356
rect 188286 465354 188292 465356
rect 78876 465294 188292 465354
rect 78876 465292 78882 465294
rect 188286 465292 188292 465294
rect 188356 465292 188362 465356
rect 91185 465220 91251 465221
rect 91134 465218 91140 465220
rect 91094 465158 91140 465218
rect 91204 465216 91251 465220
rect 91246 465160 91251 465216
rect 91134 465156 91140 465158
rect 91204 465156 91251 465160
rect 93526 465156 93532 465220
rect 93596 465218 93602 465220
rect 93669 465218 93735 465221
rect 96153 465220 96219 465221
rect 101305 465220 101371 465221
rect 103697 465220 103763 465221
rect 96102 465218 96108 465220
rect 93596 465216 93735 465218
rect 93596 465160 93674 465216
rect 93730 465160 93735 465216
rect 93596 465158 93735 465160
rect 96062 465158 96108 465218
rect 96172 465216 96219 465220
rect 101254 465218 101260 465220
rect 96214 465160 96219 465216
rect 93596 465156 93602 465158
rect 91185 465155 91251 465156
rect 93669 465155 93735 465158
rect 96102 465156 96108 465158
rect 96172 465156 96219 465160
rect 101214 465158 101260 465218
rect 101324 465216 101371 465220
rect 103646 465218 103652 465220
rect 101366 465160 101371 465216
rect 101254 465156 101260 465158
rect 101324 465156 101371 465160
rect 103606 465158 103652 465218
rect 103716 465216 103763 465220
rect 103758 465160 103763 465216
rect 103646 465156 103652 465158
rect 103716 465156 103763 465160
rect 96153 465155 96219 465156
rect 101305 465155 101371 465156
rect 103697 465155 103763 465156
rect 106181 465220 106247 465221
rect 108481 465220 108547 465221
rect 111057 465220 111123 465221
rect 128721 465220 128787 465221
rect 136081 465220 136147 465221
rect 141049 465220 141115 465221
rect 146017 465220 146083 465221
rect 106181 465216 106228 465220
rect 106292 465218 106298 465220
rect 108430 465218 108436 465220
rect 106181 465160 106186 465216
rect 106181 465156 106228 465160
rect 106292 465158 106338 465218
rect 108390 465158 108436 465218
rect 108500 465216 108547 465220
rect 111006 465218 111012 465220
rect 108542 465160 108547 465216
rect 106292 465156 106298 465158
rect 108430 465156 108436 465158
rect 108500 465156 108547 465160
rect 110966 465158 111012 465218
rect 111076 465216 111123 465220
rect 128670 465218 128676 465220
rect 111118 465160 111123 465216
rect 111006 465156 111012 465158
rect 111076 465156 111123 465160
rect 128630 465158 128676 465218
rect 128740 465216 128787 465220
rect 136030 465218 136036 465220
rect 128782 465160 128787 465216
rect 128670 465156 128676 465158
rect 128740 465156 128787 465160
rect 135990 465158 136036 465218
rect 136100 465216 136147 465220
rect 140998 465218 141004 465220
rect 136142 465160 136147 465216
rect 136030 465156 136036 465158
rect 136100 465156 136147 465160
rect 140958 465158 141004 465218
rect 141068 465216 141115 465220
rect 145966 465218 145972 465220
rect 141110 465160 141115 465216
rect 140998 465156 141004 465158
rect 141068 465156 141115 465160
rect 145926 465158 145972 465218
rect 146036 465216 146083 465220
rect 146078 465160 146083 465216
rect 145966 465156 145972 465158
rect 146036 465156 146083 465160
rect 153326 465156 153332 465220
rect 153396 465218 153402 465220
rect 154481 465218 154547 465221
rect 168465 465220 168531 465221
rect 169753 465220 169819 465221
rect 168414 465218 168420 465220
rect 153396 465216 154547 465218
rect 153396 465160 154486 465216
rect 154542 465160 154547 465216
rect 153396 465158 154547 465160
rect 168374 465158 168420 465218
rect 168484 465216 168531 465220
rect 169702 465218 169708 465220
rect 168526 465160 168531 465216
rect 153396 465156 153402 465158
rect 106181 465155 106247 465156
rect 108481 465155 108547 465156
rect 111057 465155 111123 465156
rect 128721 465155 128787 465156
rect 136081 465155 136147 465156
rect 141049 465155 141115 465156
rect 146017 465155 146083 465156
rect 154481 465155 154547 465158
rect 168414 465156 168420 465158
rect 168484 465156 168531 465160
rect 169662 465158 169708 465218
rect 169772 465216 169819 465220
rect 169814 465160 169819 465216
rect 169702 465156 169708 465158
rect 169772 465156 169819 465160
rect 180926 465156 180932 465220
rect 180996 465218 181002 465220
rect 187734 465218 187740 465220
rect 180996 465158 187740 465218
rect 180996 465156 181002 465158
rect 187734 465156 187740 465158
rect 187804 465156 187810 465220
rect 168465 465155 168531 465156
rect 169753 465155 169819 465156
rect 237373 464810 237439 464813
rect 237373 464808 240242 464810
rect 237373 464752 237378 464808
rect 237434 464752 240242 464808
rect 237373 464750 240242 464752
rect 237373 464747 237439 464750
rect 240182 464168 240242 464750
rect 131113 463996 131179 463997
rect 131062 463994 131068 463996
rect 131022 463934 131068 463994
rect 131132 463992 131179 463996
rect 131174 463936 131179 463992
rect 131062 463932 131068 463934
rect 131132 463932 131179 463936
rect 131113 463931 131179 463932
rect 83457 463724 83523 463725
rect 88517 463724 88583 463725
rect 83456 463660 83462 463724
rect 83526 463722 83532 463724
rect 88488 463722 88494 463724
rect 83526 463662 83614 463722
rect 88426 463662 88494 463722
rect 88558 463720 88583 463724
rect 88578 463664 88583 463720
rect 83526 463660 83532 463662
rect 88488 463660 88494 463662
rect 88558 463660 88583 463664
rect 83457 463659 83523 463660
rect 88517 463659 88583 463660
rect 98545 463724 98611 463725
rect 113633 463724 113699 463725
rect 116117 463724 116183 463725
rect 118601 463724 118667 463725
rect 120993 463724 121059 463725
rect 123569 463724 123635 463725
rect 125961 463724 126027 463725
rect 133505 463724 133571 463725
rect 138473 463724 138539 463725
rect 143625 463724 143691 463725
rect 148501 463724 148567 463725
rect 98545 463720 98558 463724
rect 98622 463722 98628 463724
rect 98545 463664 98550 463720
rect 98545 463660 98558 463664
rect 98622 463662 98702 463722
rect 113633 463720 113654 463724
rect 113718 463722 113724 463724
rect 116096 463722 116102 463724
rect 113633 463664 113638 463720
rect 98622 463660 98628 463662
rect 113633 463660 113654 463664
rect 113718 463662 113790 463722
rect 116026 463662 116102 463722
rect 116166 463720 116183 463724
rect 118544 463722 118550 463724
rect 116178 463664 116183 463720
rect 113718 463660 113724 463662
rect 116096 463660 116102 463662
rect 116166 463660 116183 463664
rect 118510 463662 118550 463722
rect 118614 463720 118667 463724
rect 118662 463664 118667 463720
rect 118544 463660 118550 463662
rect 118614 463660 118667 463664
rect 120992 463660 120998 463724
rect 121062 463722 121068 463724
rect 121062 463662 121150 463722
rect 123569 463720 123582 463724
rect 123646 463722 123652 463724
rect 125888 463722 125894 463724
rect 123569 463664 123574 463720
rect 121062 463660 121068 463662
rect 123569 463660 123582 463664
rect 123646 463662 123726 463722
rect 125870 463662 125894 463722
rect 123646 463660 123652 463662
rect 125888 463660 125894 463662
rect 125958 463720 126027 463724
rect 125958 463664 125966 463720
rect 126022 463664 126027 463720
rect 125958 463660 126027 463664
rect 133504 463660 133510 463724
rect 133574 463722 133580 463724
rect 138400 463722 138406 463724
rect 133574 463662 133662 463722
rect 138382 463662 138406 463722
rect 133574 463660 133580 463662
rect 138400 463660 138406 463662
rect 138470 463720 138539 463724
rect 143568 463722 143574 463724
rect 138470 463664 138478 463720
rect 138534 463664 138539 463720
rect 138470 463660 138539 463664
rect 143534 463662 143574 463722
rect 143638 463720 143691 463724
rect 148464 463722 148470 463724
rect 143686 463664 143691 463720
rect 143568 463660 143574 463662
rect 143638 463660 143691 463664
rect 148410 463662 148470 463722
rect 148534 463720 148567 463724
rect 148562 463664 148567 463720
rect 148464 463660 148470 463662
rect 148534 463660 148567 463664
rect 98545 463659 98611 463660
rect 113633 463659 113699 463660
rect 116117 463659 116183 463660
rect 118601 463659 118667 463660
rect 120993 463659 121059 463660
rect 123569 463659 123635 463660
rect 125961 463659 126027 463660
rect 133505 463659 133571 463660
rect 138473 463659 138539 463660
rect 143625 463659 143691 463660
rect 148501 463659 148567 463660
rect -960 462634 480 462724
rect 3601 462634 3667 462637
rect -960 462632 3667 462634
rect -960 462576 3606 462632
rect 3662 462576 3667 462632
rect -960 462574 3667 462576
rect -960 462484 480 462574
rect 3601 462571 3667 462574
rect 237373 462634 237439 462637
rect 240182 462634 240242 463216
rect 237373 462632 240242 462634
rect 237373 462576 237378 462632
rect 237434 462576 240242 462632
rect 237373 462574 240242 462576
rect 237373 462571 237439 462574
rect 240182 461546 240242 462128
rect 219390 461486 240242 461546
rect 186814 460940 186820 461004
rect 186884 461002 186890 461004
rect 219390 461002 219450 461486
rect 186884 460942 219450 461002
rect 186884 460940 186890 460942
rect 237465 459506 237531 459509
rect 237465 459504 240242 459506
rect 237465 459448 237470 459504
rect 237526 459448 240242 459504
rect 237465 459446 240242 459448
rect 237465 459443 237531 459446
rect 189073 459234 189139 459237
rect 187190 459232 189139 459234
rect 187190 459220 189078 459232
rect 186588 459176 189078 459220
rect 189134 459176 189139 459232
rect 186588 459174 189139 459176
rect 186588 459160 187250 459174
rect 189073 459171 189139 459174
rect 240182 459136 240242 459446
rect 237373 458282 237439 458285
rect 237373 458280 240242 458282
rect 237373 458224 237378 458280
rect 237434 458224 240242 458280
rect 237373 458222 240242 458224
rect 237373 458219 237439 458222
rect 240182 458184 240242 458222
rect 583520 457996 584960 458236
rect 238150 456860 238156 456924
rect 238220 456922 238226 456924
rect 240182 456922 240242 457096
rect 238220 456862 240242 456922
rect 238220 456860 238226 456862
rect 238017 454746 238083 454749
rect 238017 454744 240242 454746
rect 238017 454688 238022 454744
rect 238078 454688 240242 454744
rect 238017 454686 240242 454688
rect 238017 454683 238083 454686
rect 240182 454104 240242 454686
rect 238017 452706 238083 452709
rect 240182 452706 240242 453016
rect 238017 452704 240242 452706
rect 238017 452648 238022 452704
rect 238078 452648 240242 452704
rect 238017 452646 240242 452648
rect 238017 452643 238083 452646
rect 238334 451420 238340 451484
rect 238404 451482 238410 451484
rect 240182 451482 240242 452064
rect 238404 451422 240242 451482
rect 238404 451420 238410 451422
rect -960 449578 480 449668
rect 3325 449578 3391 449581
rect -960 449576 3391 449578
rect -960 449520 3330 449576
rect 3386 449520 3391 449576
rect -960 449518 3391 449520
rect -960 449428 480 449518
rect 3325 449515 3391 449518
rect 237373 449578 237439 449581
rect 237373 449576 240242 449578
rect 237373 449520 237378 449576
rect 237434 449520 240242 449576
rect 237373 449518 240242 449520
rect 237373 449515 237439 449518
rect 240182 448936 240242 449518
rect 237373 447402 237439 447405
rect 240182 447402 240242 447984
rect 237373 447400 240242 447402
rect 237373 447344 237378 447400
rect 237434 447344 240242 447400
rect 237373 447342 240242 447344
rect 237373 447339 237439 447342
rect 238293 446450 238359 446453
rect 240182 446450 240242 447032
rect 238293 446448 240242 446450
rect 238293 446392 238298 446448
rect 238354 446392 240242 446448
rect 238293 446390 240242 446392
rect 238293 446387 238359 446390
rect 583520 444668 584960 444908
rect 237373 444274 237439 444277
rect 237373 444272 240242 444274
rect 237373 444216 237378 444272
rect 237434 444216 240242 444272
rect 237373 444214 240242 444216
rect 237373 444211 237439 444214
rect 240182 443904 240242 444214
rect 237373 442370 237439 442373
rect 240182 442370 240242 442952
rect 237373 442368 240242 442370
rect 237373 442312 237378 442368
rect 237434 442312 240242 442368
rect 237373 442310 240242 442312
rect 237373 442307 237439 442310
rect 238477 441690 238543 441693
rect 240182 441690 240242 441864
rect 238477 441688 240242 441690
rect 238477 441632 238482 441688
rect 238538 441632 240242 441688
rect 238477 441630 240242 441632
rect 238477 441627 238543 441630
rect 237373 439514 237439 439517
rect 237373 439512 240242 439514
rect 237373 439456 237378 439512
rect 237434 439456 240242 439512
rect 237373 439454 240242 439456
rect 237373 439451 237439 439454
rect 240182 438872 240242 439454
rect 237373 437610 237439 437613
rect 240182 437610 240242 437784
rect 237373 437608 240242 437610
rect 237373 437552 237378 437608
rect 237434 437552 240242 437608
rect 237373 437550 240242 437552
rect 237373 437547 237439 437550
rect -960 436508 480 436748
rect 238569 436250 238635 436253
rect 240182 436250 240242 436832
rect 238569 436248 240242 436250
rect 238569 436192 238574 436248
rect 238630 436192 240242 436248
rect 238569 436190 240242 436192
rect 238569 436187 238635 436190
rect 237925 434346 237991 434349
rect 237925 434344 240242 434346
rect 237925 434288 237930 434344
rect 237986 434288 240242 434344
rect 237925 434286 240242 434288
rect 237925 434283 237991 434286
rect 240182 433840 240242 434286
rect 237373 432170 237439 432173
rect 240182 432170 240242 432752
rect 237373 432168 240242 432170
rect 237373 432112 237378 432168
rect 237434 432112 240242 432168
rect 237373 432110 240242 432112
rect 237373 432107 237439 432110
rect 237373 431218 237439 431221
rect 240182 431218 240242 431800
rect 580717 431626 580783 431629
rect 583520 431626 584960 431716
rect 580717 431624 584960 431626
rect 580717 431568 580722 431624
rect 580778 431568 584960 431624
rect 580717 431566 584960 431568
rect 580717 431563 580783 431566
rect 583520 431476 584960 431566
rect 237373 431216 240242 431218
rect 237373 431160 237378 431216
rect 237434 431160 240242 431216
rect 237373 431158 240242 431160
rect 237373 431155 237439 431158
rect 238661 429178 238727 429181
rect 238661 429176 240242 429178
rect 238661 429120 238666 429176
rect 238722 429120 240242 429176
rect 238661 429118 240242 429120
rect 238661 429115 238727 429118
rect 240182 428672 240242 429118
rect 237465 427138 237531 427141
rect 240182 427138 240242 427720
rect 237465 427136 240242 427138
rect 237465 427080 237470 427136
rect 237526 427080 240242 427136
rect 237465 427078 240242 427080
rect 237465 427075 237531 427078
rect 237373 426730 237439 426733
rect 240182 426730 240242 426768
rect 237373 426728 240242 426730
rect 237373 426672 237378 426728
rect 237434 426672 240242 426728
rect 237373 426670 240242 426672
rect 237373 426667 237439 426670
rect -960 423452 480 423692
rect 237373 423602 237439 423605
rect 240182 423602 240242 423640
rect 237373 423600 240242 423602
rect 237373 423544 237378 423600
rect 237434 423544 240242 423600
rect 237373 423542 240242 423544
rect 237373 423539 237439 423542
rect 237373 422378 237439 422381
rect 240182 422378 240242 422688
rect 237373 422376 240242 422378
rect 237373 422320 237378 422376
rect 237434 422320 240242 422376
rect 237373 422318 240242 422320
rect 237373 422315 237439 422318
rect 238661 421018 238727 421021
rect 240182 421018 240242 421600
rect 238661 421016 240242 421018
rect 238661 420960 238666 421016
rect 238722 420960 240242 421016
rect 238661 420958 240242 420960
rect 238661 420955 238727 420958
rect 237373 419250 237439 419253
rect 237373 419248 240242 419250
rect 237373 419192 237378 419248
rect 237434 419192 240242 419248
rect 237373 419190 240242 419192
rect 237373 419187 237439 419190
rect 240182 418608 240242 419190
rect 579613 418298 579679 418301
rect 583520 418298 584960 418388
rect 579613 418296 584960 418298
rect 579613 418240 579618 418296
rect 579674 418240 584960 418296
rect 579613 418238 584960 418240
rect 579613 418235 579679 418238
rect 583520 418148 584960 418238
rect 48037 416938 48103 416941
rect 237373 416938 237439 416941
rect 240182 416938 240242 417520
rect 48037 416936 49434 416938
rect 48037 416880 48042 416936
rect 48098 416924 49434 416936
rect 237373 416936 240242 416938
rect 48098 416880 50048 416924
rect 48037 416878 50048 416880
rect 48037 416875 48103 416878
rect 49374 416864 50048 416878
rect 237373 416880 237378 416936
rect 237434 416880 240242 416936
rect 237373 416878 240242 416880
rect 237373 416875 237439 416878
rect 47945 415986 48011 415989
rect 237373 415986 237439 415989
rect 240182 415986 240242 416568
rect 47945 415984 49434 415986
rect 47945 415928 47950 415984
rect 48006 415972 49434 415984
rect 237373 415984 240242 415986
rect 48006 415928 50048 415972
rect 47945 415926 50048 415928
rect 47945 415923 48011 415926
rect 49374 415912 50048 415926
rect 237373 415928 237378 415984
rect 237434 415928 240242 415984
rect 237373 415926 240242 415928
rect 237373 415923 237439 415926
rect 237373 413946 237439 413949
rect 237373 413944 240242 413946
rect 237373 413888 237378 413944
rect 237434 413888 240242 413944
rect 237373 413886 240242 413888
rect 237373 413883 237439 413886
rect 48221 413810 48287 413813
rect 48221 413808 49434 413810
rect 48221 413752 48226 413808
rect 48282 413796 49434 413808
rect 48282 413752 50048 413796
rect 48221 413750 50048 413752
rect 48221 413747 48287 413750
rect 49374 413736 50048 413750
rect 240182 413576 240242 413886
rect 49325 412858 49391 412861
rect 49325 412856 49802 412858
rect 49325 412800 49330 412856
rect 49386 412844 49802 412856
rect 49386 412800 50048 412844
rect 49325 412798 50048 412800
rect 49325 412795 49391 412798
rect 49742 412784 50048 412798
rect 237373 411906 237439 411909
rect 240182 411906 240242 412488
rect 237373 411904 240242 411906
rect 237373 411848 237378 411904
rect 237434 411848 240242 411904
rect 237373 411846 240242 411848
rect 237373 411843 237439 411846
rect 237925 411362 237991 411365
rect 240182 411362 240242 411536
rect 237925 411360 240242 411362
rect 237925 411304 237930 411360
rect 237986 411304 240242 411360
rect 237925 411302 240242 411304
rect 237925 411299 237991 411302
rect 49417 411076 49483 411079
rect 49417 411074 50048 411076
rect 49417 411018 49422 411074
rect 49478 411018 50048 411074
rect 49417 411016 50048 411018
rect 49417 411013 49483 411016
rect -960 410546 480 410636
rect 3693 410546 3759 410549
rect -960 410544 3759 410546
rect -960 410488 3698 410544
rect 3754 410488 3759 410544
rect -960 410486 3759 410488
rect -960 410396 480 410486
rect 3693 410483 3759 410486
rect 49233 410002 49299 410005
rect 49233 410000 49802 410002
rect 49233 409944 49238 410000
rect 49294 409988 49802 410000
rect 49294 409944 50048 409988
rect 49233 409942 50048 409944
rect 49233 409939 49299 409942
rect 49742 409928 50048 409942
rect 237373 408506 237439 408509
rect 237373 408504 240242 408506
rect 237373 408448 237378 408504
rect 237434 408448 240242 408504
rect 237373 408446 240242 408448
rect 237373 408443 237439 408446
rect 240182 408408 240242 408446
rect 49601 408220 49667 408223
rect 49601 408218 50048 408220
rect 49601 408162 49606 408218
rect 49662 408162 50048 408218
rect 49601 408160 50048 408162
rect 49601 408157 49667 408160
rect 237833 407146 237899 407149
rect 240182 407146 240242 407456
rect 237833 407144 240242 407146
rect 237833 407088 237838 407144
rect 237894 407088 240242 407144
rect 237833 407086 240242 407088
rect 237833 407083 237899 407086
rect 237373 405786 237439 405789
rect 240182 405786 240242 406368
rect 237373 405784 240242 405786
rect 237373 405728 237378 405784
rect 237434 405728 240242 405784
rect 237373 405726 240242 405728
rect 237373 405723 237439 405726
rect 583520 404820 584960 405060
rect 238385 404018 238451 404021
rect 238385 404016 240242 404018
rect 238385 403960 238390 404016
rect 238446 403960 240242 404016
rect 238385 403958 240242 403960
rect 238385 403955 238451 403958
rect 240182 403376 240242 403958
rect 237373 401842 237439 401845
rect 240182 401842 240242 402424
rect 237373 401840 240242 401842
rect 237373 401784 237378 401840
rect 237434 401784 240242 401840
rect 237373 401782 240242 401784
rect 237373 401779 237439 401782
rect 237373 400754 237439 400757
rect 240182 400754 240242 401336
rect 237373 400752 240242 400754
rect 237373 400696 237378 400752
rect 237434 400696 240242 400752
rect 237373 400694 240242 400696
rect 237373 400691 237439 400694
rect 189073 399394 189139 399397
rect 187190 399392 189139 399394
rect 187190 399380 189078 399392
rect 186588 399336 189078 399380
rect 189134 399336 189139 399392
rect 186588 399334 189139 399336
rect 186588 399320 187250 399334
rect 189073 399331 189139 399334
rect 238201 398850 238267 398853
rect 238201 398848 240242 398850
rect 238201 398792 238206 398848
rect 238262 398792 240242 398848
rect 238201 398790 240242 398792
rect 238201 398787 238267 398790
rect 240182 398344 240242 398790
rect 189073 397762 189139 397765
rect 187190 397760 189139 397762
rect 187190 397748 189078 397760
rect 186588 397704 189078 397748
rect 189134 397704 189139 397760
rect 186588 397702 189139 397704
rect 186588 397688 187250 397702
rect 189073 397699 189139 397702
rect -960 397490 480 397580
rect 3325 397490 3391 397493
rect -960 397488 3391 397490
rect -960 397432 3330 397488
rect 3386 397432 3391 397488
rect -960 397430 3391 397432
rect -960 397340 480 397430
rect 3325 397427 3391 397430
rect 237465 396674 237531 396677
rect 240182 396674 240242 397256
rect 237465 396672 240242 396674
rect 237465 396616 237470 396672
rect 237526 396616 240242 396672
rect 237465 396614 240242 396616
rect 237465 396611 237531 396614
rect 189073 396402 189139 396405
rect 187190 396400 189139 396402
rect 187190 396388 189078 396400
rect 186588 396344 189078 396388
rect 189134 396344 189139 396400
rect 186588 396342 189139 396344
rect 186588 396328 187250 396342
rect 189073 396339 189139 396342
rect 237373 396266 237439 396269
rect 240182 396266 240242 396304
rect 237373 396264 240242 396266
rect 237373 396208 237378 396264
rect 237434 396208 240242 396264
rect 237373 396206 240242 396208
rect 237373 396203 237439 396206
rect 189441 394906 189507 394909
rect 187190 394904 189507 394906
rect 187190 394892 189446 394904
rect 186588 394848 189446 394892
rect 189502 394848 189507 394904
rect 186588 394846 189507 394848
rect 186588 394832 187250 394846
rect 189441 394843 189507 394846
rect 238109 393954 238175 393957
rect 238109 393952 240242 393954
rect 238109 393896 238114 393952
rect 238170 393896 240242 393952
rect 238109 393894 240242 393896
rect 238109 393891 238175 393894
rect 189073 393682 189139 393685
rect 187190 393680 189139 393682
rect 187190 393668 189078 393680
rect 186588 393624 189078 393668
rect 189134 393624 189139 393680
rect 186588 393622 189139 393624
rect 186588 393608 187250 393622
rect 189073 393619 189139 393622
rect 240182 393312 240242 393894
rect 237373 392186 237439 392189
rect 240182 392186 240242 392224
rect 237373 392184 240242 392186
rect 237373 392128 237378 392184
rect 237434 392128 240242 392184
rect 237373 392126 240242 392128
rect 237373 392123 237439 392126
rect 583520 391628 584960 391868
rect 237373 390690 237439 390693
rect 240182 390690 240242 391272
rect 237373 390688 240242 390690
rect 237373 390632 237378 390688
rect 237434 390632 240242 390688
rect 237373 390630 240242 390632
rect 237373 390627 237439 390630
rect 48129 390010 48195 390013
rect 48129 390008 49434 390010
rect 48129 389952 48134 390008
rect 48190 389996 49434 390008
rect 48190 389952 50048 389996
rect 48129 389950 50048 389952
rect 48129 389947 48195 389950
rect 49374 389936 50048 389950
rect 237373 388786 237439 388789
rect 237373 388784 240242 388786
rect 237373 388728 237378 388784
rect 237434 388728 240242 388784
rect 237373 388726 240242 388728
rect 237373 388723 237439 388726
rect 47577 388378 47643 388381
rect 47577 388376 49434 388378
rect 47577 388320 47582 388376
rect 47638 388364 49434 388376
rect 47638 388320 50048 388364
rect 47577 388318 50048 388320
rect 47577 388315 47643 388318
rect 49374 388304 50048 388318
rect 240182 388144 240242 388726
rect 47853 388106 47919 388109
rect 47853 388104 49434 388106
rect 47853 388048 47858 388104
rect 47914 388092 49434 388104
rect 47914 388048 50048 388092
rect 47853 388046 50048 388048
rect 47853 388043 47919 388046
rect 49374 388032 50048 388046
rect 237373 386610 237439 386613
rect 240182 386610 240242 387192
rect 237373 386608 240242 386610
rect 237373 386552 237378 386608
rect 237434 386552 240242 386608
rect 237373 386550 240242 386552
rect 237373 386547 237439 386550
rect 237373 385522 237439 385525
rect 240182 385522 240242 386104
rect 237373 385520 240242 385522
rect 237373 385464 237378 385520
rect 237434 385464 240242 385520
rect 237373 385462 240242 385464
rect 237373 385459 237439 385462
rect -960 384284 480 384524
rect 237373 383618 237439 383621
rect 237373 383616 240242 383618
rect 237373 383560 237378 383616
rect 237434 383560 240242 383616
rect 237373 383558 240242 383560
rect 237373 383555 237439 383558
rect 240182 383112 240242 383558
rect 237465 381578 237531 381581
rect 240182 381578 240242 382160
rect 237465 381576 240242 381578
rect 237465 381520 237470 381576
rect 237526 381520 240242 381576
rect 237465 381518 240242 381520
rect 237465 381515 237531 381518
rect 237373 381034 237439 381037
rect 240182 381034 240242 381072
rect 237373 381032 240242 381034
rect 237373 380976 237378 381032
rect 237434 380976 240242 381032
rect 237373 380974 240242 380976
rect 237373 380971 237439 380974
rect 110965 379676 111031 379677
rect 113541 379676 113607 379677
rect 118325 379676 118391 379677
rect 120993 379676 121059 379677
rect 123477 379676 123543 379677
rect 130929 379676 130995 379677
rect 110928 379674 110934 379676
rect 110874 379614 110934 379674
rect 110998 379672 111031 379676
rect 113512 379674 113518 379676
rect 111026 379616 111031 379672
rect 110928 379612 110934 379614
rect 110998 379612 111031 379616
rect 113450 379614 113518 379674
rect 113582 379672 113607 379676
rect 118272 379674 118278 379676
rect 113602 379616 113607 379672
rect 113512 379612 113518 379614
rect 113582 379612 113607 379616
rect 118234 379614 118278 379674
rect 118342 379672 118391 379676
rect 118386 379616 118391 379672
rect 118272 379612 118278 379614
rect 118342 379612 118391 379616
rect 120992 379612 120998 379676
rect 121062 379674 121068 379676
rect 123440 379674 123446 379676
rect 121062 379614 121150 379674
rect 123386 379614 123446 379674
rect 123510 379672 123543 379676
rect 130920 379674 130926 379676
rect 123538 379616 123543 379672
rect 121062 379612 121068 379614
rect 123440 379612 123446 379614
rect 123510 379612 123543 379616
rect 130838 379614 130926 379674
rect 130920 379612 130926 379614
rect 130990 379612 130996 379676
rect 143432 379612 143438 379676
rect 143502 379674 143508 379676
rect 144913 379674 144979 379677
rect 143502 379672 144979 379674
rect 143502 379616 144918 379672
rect 144974 379616 144979 379672
rect 143502 379614 144979 379616
rect 143502 379612 143508 379614
rect 110965 379611 111031 379612
rect 113541 379611 113607 379612
rect 118325 379611 118391 379612
rect 120993 379611 121059 379612
rect 123477 379611 123543 379612
rect 130929 379611 130995 379612
rect 144913 379611 144979 379614
rect 87045 379540 87111 379541
rect 88149 379540 88215 379541
rect 86992 379538 86998 379540
rect 86954 379478 86998 379538
rect 87062 379536 87111 379540
rect 88080 379538 88086 379540
rect 87106 379480 87111 379536
rect 86992 379476 86998 379478
rect 87062 379476 87111 379480
rect 88058 379478 88086 379538
rect 88080 379476 88086 379478
rect 88150 379536 88215 379540
rect 88150 379480 88154 379536
rect 88210 379480 88215 379536
rect 88150 379476 88215 379480
rect 87045 379475 87111 379476
rect 88149 379475 88215 379476
rect 89437 379540 89503 379541
rect 90725 379540 90791 379541
rect 116025 379540 116091 379541
rect 150985 379540 151051 379541
rect 89437 379536 89446 379540
rect 89510 379538 89516 379540
rect 90664 379538 90670 379540
rect 89437 379480 89442 379536
rect 89437 379476 89446 379480
rect 89510 379478 89594 379538
rect 90634 379478 90670 379538
rect 90734 379536 90791 379540
rect 115974 379538 115980 379540
rect 90786 379480 90791 379536
rect 89510 379476 89516 379478
rect 90664 379476 90670 379478
rect 90734 379476 90791 379480
rect 115934 379478 115980 379538
rect 116044 379536 116091 379540
rect 150934 379538 150940 379540
rect 116086 379480 116091 379536
rect 115974 379476 115980 379478
rect 116044 379476 116091 379480
rect 150894 379478 150940 379538
rect 151004 379536 151051 379540
rect 151046 379480 151051 379536
rect 150934 379476 150940 379478
rect 151004 379476 151051 379480
rect 89437 379475 89503 379476
rect 90725 379475 90791 379476
rect 116025 379475 116091 379476
rect 150985 379475 151051 379476
rect 101254 379340 101260 379404
rect 101324 379402 101330 379404
rect 238477 379402 238543 379405
rect 101324 379400 238543 379402
rect 101324 379344 238482 379400
rect 238538 379344 238543 379400
rect 101324 379342 238543 379344
rect 101324 379340 101330 379342
rect 238477 379339 238543 379342
rect 103278 379204 103284 379268
rect 103348 379266 103354 379268
rect 238334 379266 238340 379268
rect 103348 379206 238340 379266
rect 103348 379204 103354 379206
rect 238334 379204 238340 379206
rect 238404 379204 238410 379268
rect 109166 379068 109172 379132
rect 109236 379130 109242 379132
rect 235625 379130 235691 379133
rect 109236 379128 235691 379130
rect 109236 379072 235630 379128
rect 235686 379072 235691 379128
rect 109236 379070 235691 379072
rect 109236 379068 109242 379070
rect 235625 379067 235691 379070
rect 98678 378932 98684 378996
rect 98748 378994 98754 378996
rect 189993 378994 190059 378997
rect 98748 378992 190059 378994
rect 98748 378936 189998 378992
rect 190054 378936 190059 378992
rect 98748 378934 190059 378936
rect 98748 378932 98754 378934
rect 189993 378931 190059 378934
rect 140773 378722 140839 378725
rect 238661 378722 238727 378725
rect 140773 378720 238727 378722
rect 140773 378664 140778 378720
rect 140834 378664 238666 378720
rect 238722 378664 238727 378720
rect 140773 378662 238727 378664
rect 140773 378659 140839 378662
rect 238661 378659 238727 378662
rect 580165 378450 580231 378453
rect 583520 378450 584960 378540
rect 580165 378448 584960 378450
rect 580165 378392 580170 378448
rect 580226 378392 584960 378448
rect 580165 378390 584960 378392
rect 580165 378387 580231 378390
rect 583520 378300 584960 378390
rect 67214 378116 67220 378180
rect 67284 378116 67290 378180
rect 74206 378116 74212 378180
rect 74276 378116 74282 378180
rect 77702 378116 77708 378180
rect 77772 378116 77778 378180
rect 81198 378116 81204 378180
rect 81268 378116 81274 378180
rect 91870 378116 91876 378180
rect 91940 378116 91946 378180
rect 95918 378116 95924 378180
rect 95988 378116 95994 378180
rect 99782 378116 99788 378180
rect 99852 378116 99858 378180
rect 103646 378116 103652 378180
rect 103716 378116 103722 378180
rect 128486 378116 128492 378180
rect 128556 378116 128562 378180
rect 145966 378116 145972 378180
rect 146036 378116 146042 378180
rect 153326 378116 153332 378180
rect 153396 378116 153402 378180
rect 67222 378042 67282 378116
rect 67541 378042 67607 378045
rect 67222 378040 67607 378042
rect 67222 377984 67546 378040
rect 67602 377984 67607 378040
rect 67222 377982 67607 377984
rect 74214 378042 74274 378116
rect 74349 378042 74415 378045
rect 74214 378040 74415 378042
rect 74214 377984 74354 378040
rect 74410 377984 74415 378040
rect 74214 377982 74415 377984
rect 77710 378042 77770 378116
rect 81206 378045 81266 378116
rect 91878 378045 91938 378116
rect 78489 378042 78555 378045
rect 77710 378040 78555 378042
rect 77710 377984 78494 378040
rect 78550 377984 78555 378040
rect 77710 377982 78555 377984
rect 67541 377979 67607 377982
rect 74349 377979 74415 377982
rect 78489 377979 78555 377982
rect 81157 378040 81266 378045
rect 81157 377984 81162 378040
rect 81218 377984 81266 378040
rect 81157 377982 81266 377984
rect 81157 377979 81223 377982
rect 85798 377980 85804 378044
rect 85868 378042 85874 378044
rect 85941 378042 86007 378045
rect 85868 378040 86007 378042
rect 85868 377984 85946 378040
rect 86002 377984 86007 378040
rect 85868 377982 86007 377984
rect 91878 378040 91987 378045
rect 92841 378044 92907 378045
rect 93945 378044 94011 378045
rect 95233 378044 95299 378045
rect 92790 378042 92796 378044
rect 91878 377984 91926 378040
rect 91982 377984 91987 378040
rect 91878 377982 91987 377984
rect 92750 377982 92796 378042
rect 92860 378040 92907 378044
rect 92902 377984 92907 378040
rect 85868 377980 85874 377982
rect 85941 377979 86007 377982
rect 91921 377979 91987 377982
rect 92790 377980 92796 377982
rect 92860 377980 92907 377984
rect 93894 377980 93900 378044
rect 93964 378042 94011 378044
rect 95182 378042 95188 378044
rect 93964 378040 94056 378042
rect 94006 377984 94056 378040
rect 93964 377982 94056 377984
rect 95142 377982 95188 378042
rect 95252 378040 95299 378044
rect 95294 377984 95299 378040
rect 93964 377980 94011 377982
rect 95182 377980 95188 377982
rect 95252 377980 95299 377984
rect 95926 378042 95986 378116
rect 96521 378042 96587 378045
rect 97625 378044 97691 378045
rect 97574 378042 97580 378044
rect 95926 378040 96587 378042
rect 95926 377984 96526 378040
rect 96582 377984 96587 378040
rect 95926 377982 96587 377984
rect 97534 377982 97580 378042
rect 97644 378040 97691 378044
rect 97686 377984 97691 378040
rect 92841 377979 92907 377980
rect 93945 377979 94011 377980
rect 95233 377979 95299 377980
rect 96521 377979 96587 377982
rect 97574 377980 97580 377982
rect 97644 377980 97691 377984
rect 99790 378042 99850 378116
rect 99925 378042 99991 378045
rect 99790 378040 99991 378042
rect 99790 377984 99930 378040
rect 99986 377984 99991 378040
rect 99790 377982 99991 377984
rect 103654 378042 103714 378116
rect 128494 378045 128554 378116
rect 145974 378045 146034 378116
rect 153334 378045 153394 378116
rect 104801 378042 104867 378045
rect 106089 378044 106155 378045
rect 108481 378044 108547 378045
rect 125961 378044 126027 378045
rect 106038 378042 106044 378044
rect 103654 378040 104867 378042
rect 103654 377984 104806 378040
rect 104862 377984 104867 378040
rect 103654 377982 104867 377984
rect 105998 377982 106044 378042
rect 106108 378040 106155 378044
rect 108430 378042 108436 378044
rect 106150 377984 106155 378040
rect 97625 377979 97691 377980
rect 99925 377979 99991 377982
rect 104801 377979 104867 377982
rect 106038 377980 106044 377982
rect 106108 377980 106155 377984
rect 108390 377982 108436 378042
rect 108500 378040 108547 378044
rect 125910 378042 125916 378044
rect 108542 377984 108547 378040
rect 108430 377980 108436 377982
rect 108500 377980 108547 377984
rect 125870 377982 125916 378042
rect 125980 378040 126027 378044
rect 126022 377984 126027 378040
rect 125910 377980 125916 377982
rect 125980 377980 126027 377984
rect 128494 378040 128603 378045
rect 133505 378044 133571 378045
rect 136081 378044 136147 378045
rect 138657 378044 138723 378045
rect 133454 378042 133460 378044
rect 128494 377984 128542 378040
rect 128598 377984 128603 378040
rect 128494 377982 128603 377984
rect 133414 377982 133460 378042
rect 133524 378040 133571 378044
rect 136030 378042 136036 378044
rect 133566 377984 133571 378040
rect 106089 377979 106155 377980
rect 108481 377979 108547 377980
rect 125961 377979 126027 377980
rect 128537 377979 128603 377982
rect 133454 377980 133460 377982
rect 133524 377980 133571 377984
rect 135990 377982 136036 378042
rect 136100 378040 136147 378044
rect 138606 378042 138612 378044
rect 136142 377984 136147 378040
rect 136030 377980 136036 377982
rect 136100 377980 136147 377984
rect 138566 377982 138612 378042
rect 138676 378040 138723 378044
rect 138718 377984 138723 378040
rect 138606 377980 138612 377982
rect 138676 377980 138723 377984
rect 140998 377980 141004 378044
rect 141068 378042 141074 378044
rect 141141 378042 141207 378045
rect 141068 378040 141207 378042
rect 141068 377984 141146 378040
rect 141202 377984 141207 378040
rect 141068 377982 141207 377984
rect 145974 378040 146083 378045
rect 148593 378044 148659 378045
rect 148542 378042 148548 378044
rect 145974 377984 146022 378040
rect 146078 377984 146083 378040
rect 145974 377982 146083 377984
rect 148502 377982 148548 378042
rect 148612 378040 148659 378044
rect 148654 377984 148659 378040
rect 141068 377980 141074 377982
rect 133505 377979 133571 377980
rect 136081 377979 136147 377980
rect 138657 377979 138723 377980
rect 141141 377979 141207 377982
rect 146017 377979 146083 377982
rect 148542 377980 148548 377982
rect 148612 377980 148659 377984
rect 153334 378040 153443 378045
rect 155953 378044 156019 378045
rect 155902 378042 155908 378044
rect 153334 377984 153382 378040
rect 153438 377984 153443 378040
rect 153334 377982 153443 377984
rect 155862 377982 155908 378042
rect 155972 378040 156019 378044
rect 156014 377984 156019 378040
rect 148593 377979 148659 377980
rect 153377 377979 153443 377982
rect 155902 377980 155908 377982
rect 155972 377980 156019 377984
rect 155953 377979 156019 377980
rect 237373 378042 237439 378045
rect 240182 378042 240242 378080
rect 237373 378040 240242 378042
rect 237373 377984 237378 378040
rect 237434 377984 240242 378040
rect 237373 377982 240242 377984
rect 237373 377979 237439 377982
rect 96429 377908 96495 377909
rect 96429 377904 96476 377908
rect 96540 377906 96546 377908
rect 96429 377848 96434 377904
rect 96429 377844 96476 377848
rect 96540 377846 96586 377906
rect 96540 377844 96546 377846
rect 104382 377844 104388 377908
rect 104452 377906 104458 377908
rect 238150 377906 238156 377908
rect 104452 377846 238156 377906
rect 104452 377844 104458 377846
rect 238150 377844 238156 377846
rect 238220 377844 238226 377908
rect 96429 377843 96495 377844
rect 101070 377708 101076 377772
rect 101140 377770 101146 377772
rect 102041 377770 102107 377773
rect 101140 377768 102107 377770
rect 101140 377712 102046 377768
rect 102102 377712 102107 377768
rect 101140 377710 102107 377712
rect 101140 377708 101146 377710
rect 102041 377707 102107 377710
rect 106958 377708 106964 377772
rect 107028 377770 107034 377772
rect 235165 377770 235231 377773
rect 107028 377768 235231 377770
rect 107028 377712 235170 377768
rect 235226 377712 235231 377768
rect 107028 377710 235231 377712
rect 107028 377708 107034 377710
rect 235165 377707 235231 377710
rect 108062 377572 108068 377636
rect 108132 377634 108138 377636
rect 235809 377634 235875 377637
rect 108132 377632 235875 377634
rect 108132 377576 235814 377632
rect 235870 377576 235875 377632
rect 108132 377574 235875 377576
rect 108132 377572 108138 377574
rect 235809 377571 235875 377574
rect 105854 377436 105860 377500
rect 105924 377498 105930 377500
rect 186814 377498 186820 377500
rect 105924 377438 186820 377498
rect 105924 377436 105930 377438
rect 186814 377436 186820 377438
rect 186884 377436 186890 377500
rect 180701 377362 180767 377365
rect 187734 377362 187740 377364
rect 180701 377360 187740 377362
rect 180701 377304 180706 377360
rect 180762 377304 187740 377360
rect 180701 377302 187740 377304
rect 180701 377299 180767 377302
rect 187734 377300 187740 377302
rect 187804 377300 187810 377364
rect 173198 377164 173204 377228
rect 173268 377226 173274 377228
rect 173801 377226 173867 377229
rect 173268 377224 173867 377226
rect 173268 377168 173806 377224
rect 173862 377168 173867 377224
rect 173268 377166 173867 377168
rect 173268 377164 173274 377166
rect 173801 377163 173867 377166
rect 237373 377226 237439 377229
rect 237373 377224 240242 377226
rect 237373 377168 237378 377224
rect 237434 377168 240242 377224
rect 237373 377166 240242 377168
rect 237373 377163 237439 377166
rect 66161 377092 66227 377093
rect 66110 377090 66116 377092
rect 66070 377030 66116 377090
rect 66180 377088 66227 377092
rect 66222 377032 66227 377088
rect 66110 377028 66116 377030
rect 66180 377028 66227 377032
rect 68318 377028 68324 377092
rect 68388 377090 68394 377092
rect 68921 377090 68987 377093
rect 68388 377088 68987 377090
rect 68388 377032 68926 377088
rect 68982 377032 68987 377088
rect 68388 377030 68987 377032
rect 68388 377028 68394 377030
rect 66161 377027 66227 377028
rect 68921 377027 68987 377030
rect 69606 377028 69612 377092
rect 69676 377090 69682 377092
rect 70301 377090 70367 377093
rect 69676 377088 70367 377090
rect 69676 377032 70306 377088
rect 70362 377032 70367 377088
rect 69676 377030 70367 377032
rect 69676 377028 69682 377030
rect 70301 377027 70367 377030
rect 70526 377028 70532 377092
rect 70596 377090 70602 377092
rect 71681 377090 71747 377093
rect 70596 377088 71747 377090
rect 70596 377032 71686 377088
rect 71742 377032 71747 377088
rect 70596 377030 71747 377032
rect 70596 377028 70602 377030
rect 71681 377027 71747 377030
rect 71814 377028 71820 377092
rect 71884 377090 71890 377092
rect 73061 377090 73127 377093
rect 71884 377088 73127 377090
rect 71884 377032 73066 377088
rect 73122 377032 73127 377088
rect 71884 377030 73127 377032
rect 71884 377028 71890 377030
rect 73061 377027 73127 377030
rect 75494 377028 75500 377092
rect 75564 377090 75570 377092
rect 75821 377090 75887 377093
rect 75564 377088 75887 377090
rect 75564 377032 75826 377088
rect 75882 377032 75887 377088
rect 75564 377030 75887 377032
rect 75564 377028 75570 377030
rect 75821 377027 75887 377030
rect 76598 377028 76604 377092
rect 76668 377090 76674 377092
rect 77201 377090 77267 377093
rect 78305 377092 78371 377093
rect 78254 377090 78260 377092
rect 76668 377088 77267 377090
rect 76668 377032 77206 377088
rect 77262 377032 77267 377088
rect 76668 377030 77267 377032
rect 78214 377030 78260 377090
rect 78324 377088 78371 377092
rect 78366 377032 78371 377088
rect 76668 377028 76674 377030
rect 77201 377027 77267 377030
rect 78254 377028 78260 377030
rect 78324 377028 78371 377032
rect 78806 377028 78812 377092
rect 78876 377090 78882 377092
rect 79961 377090 80027 377093
rect 78876 377088 80027 377090
rect 78876 377032 79966 377088
rect 80022 377032 80027 377088
rect 78876 377030 80027 377032
rect 78876 377028 78882 377030
rect 78305 377027 78371 377028
rect 79961 377027 80027 377030
rect 80094 377028 80100 377092
rect 80164 377090 80170 377092
rect 81249 377090 81315 377093
rect 80164 377088 81315 377090
rect 80164 377032 81254 377088
rect 81310 377032 81315 377088
rect 80164 377030 81315 377032
rect 80164 377028 80170 377030
rect 81249 377027 81315 377030
rect 82486 377028 82492 377092
rect 82556 377090 82562 377092
rect 82721 377090 82787 377093
rect 82556 377088 82787 377090
rect 82556 377032 82726 377088
rect 82782 377032 82787 377088
rect 82556 377030 82787 377032
rect 82556 377028 82562 377030
rect 82721 377027 82787 377030
rect 83590 377028 83596 377092
rect 83660 377090 83666 377092
rect 84101 377090 84167 377093
rect 83660 377088 84167 377090
rect 83660 377032 84106 377088
rect 84162 377032 84167 377088
rect 83660 377030 84167 377032
rect 83660 377028 83666 377030
rect 84101 377027 84167 377030
rect 84510 377028 84516 377092
rect 84580 377090 84586 377092
rect 85481 377090 85547 377093
rect 84580 377088 85547 377090
rect 84580 377032 85486 377088
rect 85542 377032 85547 377088
rect 84580 377030 85547 377032
rect 84580 377028 84586 377030
rect 85481 377027 85547 377030
rect 85982 377028 85988 377092
rect 86052 377090 86058 377092
rect 86769 377090 86835 377093
rect 86052 377088 86835 377090
rect 86052 377032 86774 377088
rect 86830 377032 86835 377088
rect 86052 377030 86835 377032
rect 86052 377028 86058 377030
rect 86769 377027 86835 377030
rect 88558 377028 88564 377092
rect 88628 377090 88634 377092
rect 89621 377090 89687 377093
rect 88628 377088 89687 377090
rect 88628 377032 89626 377088
rect 89682 377032 89687 377088
rect 88628 377030 89687 377032
rect 88628 377028 88634 377030
rect 89621 377027 89687 377030
rect 91134 377028 91140 377092
rect 91204 377090 91210 377092
rect 92381 377090 92447 377093
rect 91204 377088 92447 377090
rect 91204 377032 92386 377088
rect 92442 377032 92447 377088
rect 91204 377030 92447 377032
rect 91204 377028 91210 377030
rect 92381 377027 92447 377030
rect 93526 377028 93532 377092
rect 93596 377090 93602 377092
rect 93761 377090 93827 377093
rect 93596 377088 93827 377090
rect 93596 377032 93766 377088
rect 93822 377032 93827 377088
rect 93596 377030 93827 377032
rect 93596 377028 93602 377030
rect 93761 377027 93827 377030
rect 98310 377028 98316 377092
rect 98380 377090 98386 377092
rect 99281 377090 99347 377093
rect 98380 377088 99347 377090
rect 98380 377032 99286 377088
rect 99342 377032 99347 377088
rect 98380 377030 99347 377032
rect 98380 377028 98386 377030
rect 99281 377027 99347 377030
rect 102174 377028 102180 377092
rect 102244 377090 102250 377092
rect 238293 377090 238359 377093
rect 102244 377088 238359 377090
rect 102244 377032 238298 377088
rect 238354 377032 238359 377088
rect 102244 377030 238359 377032
rect 102244 377028 102250 377030
rect 238293 377027 238359 377030
rect 240182 376992 240242 377166
rect 73102 376892 73108 376956
rect 73172 376954 73178 376956
rect 74441 376954 74507 376957
rect 73172 376952 74507 376954
rect 73172 376896 74446 376952
rect 74502 376896 74507 376952
rect 73172 376894 74507 376896
rect 73172 376892 73178 376894
rect 74441 376891 74507 376894
rect 80830 376892 80836 376956
rect 80900 376954 80906 376956
rect 81341 376954 81407 376957
rect 80900 376952 81407 376954
rect 80900 376896 81346 376952
rect 81402 376896 81407 376952
rect 80900 376894 81407 376896
rect 80900 376892 80906 376894
rect 81341 376891 81407 376894
rect 83406 376892 83412 376956
rect 83476 376954 83482 376956
rect 84009 376954 84075 376957
rect 83476 376952 84075 376954
rect 83476 376896 84014 376952
rect 84070 376896 84075 376952
rect 83476 376894 84075 376896
rect 83476 376892 83482 376894
rect 84009 376891 84075 376894
rect 173382 376892 173388 376956
rect 173452 376954 173458 376956
rect 173709 376954 173775 376957
rect 173452 376952 173775 376954
rect 173452 376896 173714 376952
rect 173770 376896 173775 376952
rect 173452 376894 173775 376896
rect 173452 376892 173458 376894
rect 173709 376891 173775 376894
rect 237373 376682 237439 376685
rect 237373 376680 240242 376682
rect 237373 376624 237378 376680
rect 237434 376624 240242 376680
rect 237373 376622 240242 376624
rect 237373 376619 237439 376622
rect 240182 376040 240242 376622
rect 237373 373690 237439 373693
rect 237373 373688 240242 373690
rect 237373 373632 237378 373688
rect 237434 373632 240242 373688
rect 237373 373630 240242 373632
rect 237373 373627 237439 373630
rect 240182 373048 240242 373630
rect 237373 372466 237439 372469
rect 237373 372464 240242 372466
rect 237373 372408 237378 372464
rect 237434 372408 240242 372464
rect 237373 372406 240242 372408
rect 237373 372403 237439 372406
rect 240182 371960 240242 372406
rect -960 371228 480 371468
rect 237373 371106 237439 371109
rect 237373 371104 240242 371106
rect 237373 371048 237378 371104
rect 237434 371048 240242 371104
rect 237373 371046 240242 371048
rect 237373 371043 237439 371046
rect 240182 371008 240242 371046
rect 237373 368386 237439 368389
rect 237373 368384 240242 368386
rect 237373 368328 237378 368384
rect 237434 368328 240242 368384
rect 237373 368326 240242 368328
rect 237373 368323 237439 368326
rect 240182 367880 240242 368326
rect 237373 367026 237439 367029
rect 237373 367024 240242 367026
rect 237373 366968 237378 367024
rect 237434 366968 240242 367024
rect 237373 366966 240242 366968
rect 237373 366963 237439 366966
rect 240182 366928 240242 366966
rect 237465 366482 237531 366485
rect 237465 366480 240242 366482
rect 237465 366424 237470 366480
rect 237526 366424 240242 366480
rect 237465 366422 240242 366424
rect 237465 366419 237531 366422
rect 240182 365840 240242 366422
rect 580165 365122 580231 365125
rect 583520 365122 584960 365212
rect 580165 365120 584960 365122
rect 580165 365064 580170 365120
rect 580226 365064 584960 365120
rect 580165 365062 584960 365064
rect 580165 365059 580231 365062
rect 583520 364972 584960 365062
rect 237373 362810 237439 362813
rect 240182 362810 240242 362848
rect 237373 362808 240242 362810
rect 237373 362752 237378 362808
rect 237434 362752 240242 362808
rect 237373 362750 240242 362752
rect 237373 362747 237439 362750
rect 237465 362538 237531 362541
rect 237465 362536 240242 362538
rect 237465 362480 237470 362536
rect 237526 362480 240242 362536
rect 237465 362478 240242 362480
rect 237465 362475 237531 362478
rect 240182 361896 240242 362478
rect 237373 361450 237439 361453
rect 237373 361448 240242 361450
rect 237373 361392 237378 361448
rect 237434 361392 240242 361448
rect 237373 361390 240242 361392
rect 237373 361387 237439 361390
rect 240182 360808 240242 361390
rect 237373 360090 237439 360093
rect 237373 360088 240242 360090
rect 237373 360032 237378 360088
rect 237434 360032 240242 360088
rect 237373 360030 240242 360032
rect 237373 360027 237439 360030
rect 240182 359856 240242 360030
rect 237373 358730 237439 358733
rect 240182 358730 240242 358768
rect 237373 358728 240242 358730
rect 237373 358672 237378 358728
rect 237434 358672 240242 358728
rect 237373 358670 240242 358672
rect 237373 358667 237439 358670
rect -960 358458 480 358548
rect 3785 358458 3851 358461
rect -960 358456 3851 358458
rect -960 358400 3790 358456
rect 3846 358400 3851 358456
rect -960 358398 3851 358400
rect -960 358308 480 358398
rect 3785 358395 3851 358398
rect 237465 358458 237531 358461
rect 237465 358456 240242 358458
rect 237465 358400 237470 358456
rect 237526 358400 240242 358456
rect 237465 358398 240242 358400
rect 237465 358395 237531 358398
rect 240182 357816 240242 358398
rect 237373 357370 237439 357373
rect 237373 357368 240242 357370
rect 237373 357312 237378 357368
rect 237434 357312 240242 357368
rect 237373 357310 240242 357312
rect 237373 357307 237439 357310
rect 240182 356728 240242 357310
rect 237373 355874 237439 355877
rect 237373 355872 240242 355874
rect 237373 355816 237378 355872
rect 237434 355816 240242 355872
rect 237373 355814 240242 355816
rect 237373 355811 237439 355814
rect 240182 355776 240242 355814
rect 237465 355330 237531 355333
rect 237465 355328 240242 355330
rect 237465 355272 237470 355328
rect 237526 355272 240242 355328
rect 237465 355270 240242 355272
rect 237465 355267 237531 355270
rect 240182 354688 240242 355270
rect 237373 354378 237439 354381
rect 237373 354376 240242 354378
rect 237373 354320 237378 354376
rect 237434 354320 240242 354376
rect 237373 354318 240242 354320
rect 237373 354315 237439 354318
rect 240182 353736 240242 354318
rect 237373 353018 237439 353021
rect 237373 353016 240242 353018
rect 237373 352960 237378 353016
rect 237434 352960 240242 353016
rect 237373 352958 240242 352960
rect 237373 352955 237439 352958
rect 240182 352648 240242 352958
rect 237373 351794 237439 351797
rect 237373 351792 240242 351794
rect 237373 351736 237378 351792
rect 237434 351736 240242 351792
rect 583520 351780 584960 352020
rect 237373 351734 240242 351736
rect 237373 351731 237439 351734
rect 240182 351696 240242 351734
rect 237465 351386 237531 351389
rect 237465 351384 240242 351386
rect 237465 351328 237470 351384
rect 237526 351328 240242 351384
rect 237465 351326 240242 351328
rect 237465 351323 237531 351326
rect 240182 350744 240242 351326
rect 237373 350298 237439 350301
rect 237373 350296 240242 350298
rect 237373 350240 237378 350296
rect 237434 350240 240242 350296
rect 237373 350238 240242 350240
rect 237373 350235 237439 350238
rect 240182 349656 240242 350238
rect 237373 349074 237439 349077
rect 237373 349072 240242 349074
rect 237373 349016 237378 349072
rect 237434 349016 240242 349072
rect 237373 349014 240242 349016
rect 237373 349011 237439 349014
rect 240182 348704 240242 349014
rect 237465 347714 237531 347717
rect 237465 347712 240242 347714
rect 237465 347656 237470 347712
rect 237526 347656 240242 347712
rect 237465 347654 240242 347656
rect 237465 347651 237531 347654
rect 240182 347616 240242 347654
rect 237373 347306 237439 347309
rect 237373 347304 240242 347306
rect 237373 347248 237378 347304
rect 237434 347248 240242 347304
rect 237373 347246 240242 347248
rect 237373 347243 237439 347246
rect 240182 346664 240242 347246
rect 237373 346218 237439 346221
rect 237373 346216 240242 346218
rect 237373 346160 237378 346216
rect 237434 346160 240242 346216
rect 237373 346158 240242 346160
rect 237373 346155 237439 346158
rect 240182 345576 240242 346158
rect -960 345402 480 345492
rect 3049 345402 3115 345405
rect -960 345400 3115 345402
rect -960 345344 3054 345400
rect 3110 345344 3115 345400
rect -960 345342 3115 345344
rect -960 345252 480 345342
rect 3049 345339 3115 345342
rect 237373 344858 237439 344861
rect 237373 344856 240242 344858
rect 237373 344800 237378 344856
rect 237434 344800 240242 344856
rect 237373 344798 240242 344800
rect 237373 344795 237439 344798
rect 240182 344624 240242 344798
rect 238017 343634 238083 343637
rect 238017 343632 240242 343634
rect 238017 343576 238022 343632
rect 238078 343576 240242 343632
rect 238017 343574 240242 343576
rect 238017 343571 238083 343574
rect 240182 343536 240242 343574
rect 237373 343226 237439 343229
rect 237373 343224 240242 343226
rect 237373 343168 237378 343224
rect 237434 343168 240242 343224
rect 237373 343166 240242 343168
rect 237373 343163 237439 343166
rect 240182 342584 240242 343166
rect 237373 342138 237439 342141
rect 237373 342136 240242 342138
rect 237373 342080 237378 342136
rect 237434 342080 240242 342136
rect 237373 342078 240242 342080
rect 237373 342075 237439 342078
rect 240182 341496 240242 342078
rect 237373 340778 237439 340781
rect 237373 340776 240242 340778
rect 237373 340720 237378 340776
rect 237434 340720 240242 340776
rect 237373 340718 240242 340720
rect 237373 340715 237439 340718
rect 240182 340544 240242 340718
rect 237465 340234 237531 340237
rect 237465 340232 240242 340234
rect 237465 340176 237470 340232
rect 237526 340176 240242 340232
rect 237465 340174 240242 340176
rect 237465 340171 237531 340174
rect 240182 339592 240242 340174
rect 238109 339146 238175 339149
rect 238109 339144 240242 339146
rect 238109 339088 238114 339144
rect 238170 339088 240242 339144
rect 238109 339086 240242 339088
rect 238109 339083 238175 339086
rect 240182 338504 240242 339086
rect 583520 338452 584960 338692
rect 237373 338058 237439 338061
rect 237373 338056 240242 338058
rect 237373 338000 237378 338056
rect 237434 338000 240242 338056
rect 237373 337998 240242 338000
rect 237373 337995 237439 337998
rect 240182 337552 240242 337998
rect 237373 336562 237439 336565
rect 237373 336560 240242 336562
rect 237373 336504 237378 336560
rect 237434 336504 240242 336560
rect 237373 336502 240242 336504
rect 237373 336499 237439 336502
rect 240182 336464 240242 336502
rect 237465 336154 237531 336157
rect 237465 336152 240242 336154
rect 237465 336096 237470 336152
rect 237526 336096 240242 336152
rect 237465 336094 240242 336096
rect 237465 336091 237531 336094
rect 240182 335512 240242 336094
rect 237373 335066 237439 335069
rect 237373 335064 240242 335066
rect 237373 335008 237378 335064
rect 237434 335008 240242 335064
rect 237373 335006 240242 335008
rect 237373 335003 237439 335006
rect 240182 334424 240242 335006
rect 237373 333842 237439 333845
rect 237373 333840 240242 333842
rect 237373 333784 237378 333840
rect 237434 333784 240242 333840
rect 237373 333782 240242 333784
rect 237373 333779 237439 333782
rect 240182 333472 240242 333782
rect 237373 332482 237439 332485
rect 237373 332480 240242 332482
rect -960 332196 480 332436
rect 237373 332424 237378 332480
rect 237434 332424 240242 332480
rect 237373 332422 240242 332424
rect 237373 332419 237439 332422
rect 240182 332384 240242 332422
rect 237465 332074 237531 332077
rect 237465 332072 240242 332074
rect 237465 332016 237470 332072
rect 237526 332016 240242 332072
rect 237465 332014 240242 332016
rect 237465 332011 237531 332014
rect 240182 331432 240242 332014
rect 237373 331122 237439 331125
rect 237373 331120 240242 331122
rect 237373 331064 237378 331120
rect 237434 331064 240242 331120
rect 237373 331062 240242 331064
rect 237373 331059 237439 331062
rect 240182 330480 240242 331062
rect 237373 329626 237439 329629
rect 237373 329624 240242 329626
rect 237373 329568 237378 329624
rect 237434 329568 240242 329624
rect 237373 329566 240242 329568
rect 237373 329563 237439 329566
rect 240182 329392 240242 329566
rect 237465 329082 237531 329085
rect 237465 329080 240242 329082
rect 237465 329024 237470 329080
rect 237526 329024 240242 329080
rect 237465 329022 240242 329024
rect 237465 329019 237531 329022
rect 240182 328440 240242 329022
rect 237373 327994 237439 327997
rect 237373 327992 240242 327994
rect 237373 327936 237378 327992
rect 237434 327936 240242 327992
rect 237373 327934 240242 327936
rect 237373 327931 237439 327934
rect 240182 327352 240242 327934
rect 237373 327042 237439 327045
rect 237373 327040 240242 327042
rect 237373 326984 237378 327040
rect 237434 326984 240242 327040
rect 237373 326982 240242 326984
rect 237373 326979 237439 326982
rect 240182 326400 240242 326982
rect 237373 325546 237439 325549
rect 237373 325544 240242 325546
rect 237373 325488 237378 325544
rect 237434 325488 240242 325544
rect 237373 325486 240242 325488
rect 237373 325483 237439 325486
rect 240182 325312 240242 325486
rect 579613 325274 579679 325277
rect 583520 325274 584960 325364
rect 579613 325272 584960 325274
rect 579613 325216 579618 325272
rect 579674 325216 584960 325272
rect 579613 325214 584960 325216
rect 579613 325211 579679 325214
rect 583520 325124 584960 325214
rect 237373 325002 237439 325005
rect 237373 325000 240242 325002
rect 237373 324944 237378 325000
rect 237434 324944 240242 325000
rect 237373 324942 240242 324944
rect 237373 324939 237439 324942
rect 240182 324360 240242 324942
rect 237373 323914 237439 323917
rect 237373 323912 240242 323914
rect 237373 323856 237378 323912
rect 237434 323856 240242 323912
rect 237373 323854 240242 323856
rect 237373 323851 237439 323854
rect 240182 323272 240242 323854
rect 237465 322826 237531 322829
rect 237465 322824 240242 322826
rect 237465 322768 237470 322824
rect 237526 322768 240242 322824
rect 237465 322766 240242 322768
rect 237465 322763 237531 322766
rect 240182 322320 240242 322766
rect 237373 321466 237439 321469
rect 237373 321464 240242 321466
rect 237373 321408 237378 321464
rect 237434 321408 240242 321464
rect 237373 321406 240242 321408
rect 237373 321403 237439 321406
rect 240182 321232 240242 321406
rect 237465 320922 237531 320925
rect 237465 320920 240242 320922
rect 237465 320864 237470 320920
rect 237526 320864 240242 320920
rect 237465 320862 240242 320864
rect 237465 320859 237531 320862
rect 240182 320280 240242 320862
rect 237373 319970 237439 319973
rect 237373 319968 240242 319970
rect 237373 319912 237378 319968
rect 237434 319912 240242 319968
rect 237373 319910 240242 319912
rect 237373 319907 237439 319910
rect -960 319140 480 319380
rect 240182 319328 240242 319910
rect 188286 317460 188292 317524
rect 188356 317522 188362 317524
rect 240182 317522 240242 318240
rect 188356 317462 240242 317522
rect 188356 317460 188362 317462
rect 237373 317386 237439 317389
rect 237373 317384 240242 317386
rect 237373 317328 237378 317384
rect 237434 317328 240242 317384
rect 237373 317326 240242 317328
rect 237373 317323 237439 317326
rect 240182 317288 240242 317326
rect 237557 316842 237623 316845
rect 237557 316840 240242 316842
rect 237557 316784 237562 316840
rect 237618 316784 240242 316840
rect 237557 316782 240242 316784
rect 237557 316779 237623 316782
rect 240182 316200 240242 316782
rect 237373 315890 237439 315893
rect 237373 315888 240242 315890
rect 237373 315832 237378 315888
rect 237434 315832 240242 315888
rect 237373 315830 240242 315832
rect 237373 315827 237439 315830
rect 240182 315248 240242 315830
rect 237373 314530 237439 314533
rect 237373 314528 240242 314530
rect 237373 314472 237378 314528
rect 237434 314472 240242 314528
rect 237373 314470 240242 314472
rect 237373 314467 237439 314470
rect 240182 314160 240242 314470
rect 237373 313170 237439 313173
rect 240182 313170 240242 313208
rect 237373 313168 240242 313170
rect 237373 313112 237378 313168
rect 237434 313112 240242 313168
rect 237373 313110 240242 313112
rect 237373 313107 237439 313110
rect 237465 312762 237531 312765
rect 237465 312760 240242 312762
rect 237465 312704 237470 312760
rect 237526 312704 240242 312760
rect 237465 312702 240242 312704
rect 237465 312699 237531 312702
rect 240182 312120 240242 312702
rect 580809 312082 580875 312085
rect 583520 312082 584960 312172
rect 580809 312080 584960 312082
rect 580809 312024 580814 312080
rect 580870 312024 584960 312080
rect 580809 312022 584960 312024
rect 580809 312019 580875 312022
rect 583520 311932 584960 312022
rect 237373 311810 237439 311813
rect 237373 311808 240242 311810
rect 237373 311752 237378 311808
rect 237434 311752 240242 311808
rect 237373 311750 240242 311752
rect 237373 311747 237439 311750
rect 240182 311168 240242 311750
rect 237373 309498 237439 309501
rect 240182 309498 240242 310080
rect 237373 309496 240242 309498
rect 237373 309440 237378 309496
rect 237434 309440 240242 309496
rect 237373 309438 240242 309440
rect 237373 309435 237439 309438
rect 237465 309226 237531 309229
rect 237465 309224 240242 309226
rect 237465 309168 237470 309224
rect 237526 309168 240242 309224
rect 237465 309166 240242 309168
rect 237465 309163 237531 309166
rect 240182 309128 240242 309166
rect 237373 307866 237439 307869
rect 240182 307866 240242 308176
rect 237373 307864 240242 307866
rect 237373 307808 237378 307864
rect 237434 307808 240242 307864
rect 237373 307806 240242 307808
rect 237373 307803 237439 307806
rect 238017 306506 238083 306509
rect 240182 306506 240242 307088
rect 238017 306504 240242 306506
rect 238017 306448 238022 306504
rect 238078 306448 240242 306504
rect 238017 306446 240242 306448
rect 238017 306443 238083 306446
rect -960 306234 480 306324
rect 3877 306234 3943 306237
rect -960 306232 3943 306234
rect -960 306176 3882 306232
rect 3938 306176 3943 306232
rect -960 306174 3943 306176
rect -960 306084 480 306174
rect 3877 306171 3943 306174
rect 237465 305554 237531 305557
rect 240182 305554 240242 306136
rect 237465 305552 240242 305554
rect 237465 305496 237470 305552
rect 237526 305496 240242 305552
rect 237465 305494 240242 305496
rect 237465 305491 237531 305494
rect 237373 305010 237439 305013
rect 240182 305010 240242 305048
rect 237373 305008 240242 305010
rect 237373 304952 237378 305008
rect 237434 304952 240242 305008
rect 237373 304950 240242 304952
rect 237373 304947 237439 304950
rect 237373 303922 237439 303925
rect 240182 303922 240242 304096
rect 237373 303920 240242 303922
rect 237373 303864 237378 303920
rect 237434 303864 240242 303920
rect 237373 303862 240242 303864
rect 237373 303859 237439 303862
rect 237373 302426 237439 302429
rect 240182 302426 240242 303008
rect 237373 302424 240242 302426
rect 237373 302368 237378 302424
rect 237434 302368 240242 302424
rect 237373 302366 240242 302368
rect 237373 302363 237439 302366
rect 237465 301474 237531 301477
rect 240182 301474 240242 302056
rect 237465 301472 240242 301474
rect 237465 301416 237470 301472
rect 237526 301416 240242 301472
rect 237465 301414 240242 301416
rect 237465 301411 237531 301414
rect 237373 300930 237439 300933
rect 240182 300930 240242 300968
rect 237373 300928 240242 300930
rect 237373 300872 237378 300928
rect 237434 300872 240242 300928
rect 237373 300870 240242 300872
rect 237373 300867 237439 300870
rect 236729 300114 236795 300117
rect 236729 300112 240242 300114
rect 236729 300056 236734 300112
rect 236790 300056 240242 300112
rect 236729 300054 240242 300056
rect 236729 300051 236795 300054
rect 240182 300016 240242 300054
rect 239814 298898 240212 298958
rect 237373 298890 237439 298893
rect 239814 298890 239874 298898
rect 237373 298888 239874 298890
rect 237373 298832 237378 298888
rect 237434 298832 239874 298888
rect 237373 298830 239874 298832
rect 237373 298827 237439 298830
rect 583520 298604 584960 298844
rect 239814 297946 240212 298006
rect 237373 297938 237439 297941
rect 239814 297938 239874 297946
rect 237373 297936 239874 297938
rect 237373 297880 237378 297936
rect 237434 297880 239874 297936
rect 237373 297878 239874 297880
rect 237373 297875 237439 297878
rect 239814 296994 240212 297054
rect 236821 296986 236887 296989
rect 239814 296986 239874 296994
rect 236821 296984 239874 296986
rect 236821 296928 236826 296984
rect 236882 296928 239874 296984
rect 236821 296926 239874 296928
rect 236821 296923 236887 296926
rect 239814 295906 240212 295966
rect 237373 295898 237439 295901
rect 239814 295898 239874 295906
rect 237373 295896 239874 295898
rect 237373 295840 237378 295896
rect 237434 295840 239874 295896
rect 237373 295838 239874 295840
rect 237373 295835 237439 295838
rect 239814 294954 240212 295014
rect 237373 294946 237439 294949
rect 239814 294946 239874 294954
rect 237373 294944 239874 294946
rect 237373 294888 237378 294944
rect 237434 294888 239874 294944
rect 237373 294886 239874 294888
rect 237373 294883 237439 294886
rect 239814 293866 240212 293926
rect 236913 293858 236979 293861
rect 239814 293858 239874 293866
rect 236913 293856 239874 293858
rect 236913 293800 236918 293856
rect 236974 293800 239874 293856
rect 236913 293798 239874 293800
rect 236913 293795 236979 293798
rect -960 293178 480 293268
rect 3141 293178 3207 293181
rect -960 293176 3207 293178
rect -960 293120 3146 293176
rect 3202 293120 3207 293176
rect -960 293118 3207 293120
rect -960 293028 480 293118
rect 3141 293115 3207 293118
rect 239814 292914 240212 292974
rect 237373 292906 237439 292909
rect 239814 292906 239874 292914
rect 237373 292904 239874 292906
rect 237373 292848 237378 292904
rect 237434 292848 239874 292904
rect 237373 292846 239874 292848
rect 237373 292843 237439 292846
rect 239814 291826 240212 291886
rect 237373 291818 237439 291821
rect 239814 291818 239874 291826
rect 237373 291816 239874 291818
rect 237373 291760 237378 291816
rect 237434 291760 239874 291816
rect 237373 291758 239874 291760
rect 237373 291755 237439 291758
rect 239814 290874 240212 290934
rect 237005 290866 237071 290869
rect 239814 290866 239874 290874
rect 237005 290864 239874 290866
rect 237005 290808 237010 290864
rect 237066 290808 239874 290864
rect 237005 290806 239874 290808
rect 237005 290803 237071 290806
rect 237373 289914 237439 289917
rect 237373 289912 239874 289914
rect 237373 289856 237378 289912
rect 237434 289856 239874 289912
rect 237373 289854 239874 289856
rect 237373 289851 237439 289854
rect 239814 289846 239874 289854
rect 239814 289786 240212 289846
rect 239814 288834 240212 288894
rect 237373 288826 237439 288829
rect 239814 288826 239874 288834
rect 237373 288824 239874 288826
rect 237373 288768 237378 288824
rect 237434 288768 239874 288824
rect 237373 288766 239874 288768
rect 237373 288763 237439 288766
rect 239814 287746 240212 287806
rect 237097 287738 237163 287741
rect 239814 287738 239874 287746
rect 237097 287736 239874 287738
rect 237097 287680 237102 287736
rect 237158 287680 239874 287736
rect 237097 287678 239874 287680
rect 237097 287675 237163 287678
rect 239814 286794 240212 286854
rect 237465 286786 237531 286789
rect 239814 286786 239874 286794
rect 237465 286784 239874 286786
rect 237465 286728 237470 286784
rect 237526 286728 239874 286784
rect 237465 286726 239874 286728
rect 237465 286723 237531 286726
rect 116158 286452 116164 286516
rect 116228 286514 116234 286516
rect 117221 286514 117287 286517
rect 116228 286512 117287 286514
rect 116228 286456 117226 286512
rect 117282 286456 117287 286512
rect 116228 286454 117287 286456
rect 116228 286452 116234 286454
rect 117221 286451 117287 286454
rect 136030 286316 136036 286380
rect 136100 286378 136106 286380
rect 136541 286378 136607 286381
rect 136100 286376 136607 286378
rect 136100 286320 136546 286376
rect 136602 286320 136607 286376
rect 136100 286318 136607 286320
rect 136100 286316 136106 286318
rect 136541 286315 136607 286318
rect 169702 286316 169708 286380
rect 169772 286378 169778 286380
rect 170673 286378 170739 286381
rect 169772 286376 170739 286378
rect 169772 286320 170678 286376
rect 170734 286320 170739 286376
rect 169772 286318 170739 286320
rect 169772 286316 169778 286318
rect 170673 286315 170739 286318
rect 168414 286180 168420 286244
rect 168484 286242 168490 286244
rect 169661 286242 169727 286245
rect 168484 286240 169727 286242
rect 168484 286184 169666 286240
rect 169722 286184 169727 286240
rect 168484 286182 169727 286184
rect 168484 286180 168490 286182
rect 169661 286179 169727 286182
rect 125910 286044 125916 286108
rect 125980 286106 125986 286108
rect 126881 286106 126947 286109
rect 125980 286104 126947 286106
rect 125980 286048 126886 286104
rect 126942 286048 126947 286104
rect 125980 286046 126947 286048
rect 125980 286044 125986 286046
rect 126881 286043 126947 286046
rect 131062 286044 131068 286108
rect 131132 286106 131138 286108
rect 132309 286106 132375 286109
rect 131132 286104 132375 286106
rect 131132 286048 132314 286104
rect 132370 286048 132375 286104
rect 131132 286046 132375 286048
rect 131132 286044 131138 286046
rect 132309 286043 132375 286046
rect 133454 286044 133460 286108
rect 133524 286106 133530 286108
rect 133781 286106 133847 286109
rect 133524 286104 133847 286106
rect 133524 286048 133786 286104
rect 133842 286048 133847 286104
rect 133524 286046 133847 286048
rect 133524 286044 133530 286046
rect 133781 286043 133847 286046
rect 108430 285908 108436 285972
rect 108500 285970 108506 285972
rect 108941 285970 109007 285973
rect 108500 285968 109007 285970
rect 108500 285912 108946 285968
rect 109002 285912 109007 285968
rect 108500 285910 109007 285912
rect 108500 285908 108506 285910
rect 108941 285907 109007 285910
rect 111006 285908 111012 285972
rect 111076 285970 111082 285972
rect 111701 285970 111767 285973
rect 111076 285968 111767 285970
rect 111076 285912 111706 285968
rect 111762 285912 111767 285968
rect 111076 285910 111767 285912
rect 111076 285908 111082 285910
rect 111701 285907 111767 285910
rect 237373 285970 237439 285973
rect 237373 285968 239874 285970
rect 237373 285912 237378 285968
rect 237434 285912 239874 285968
rect 237373 285910 239874 285912
rect 237373 285907 237439 285910
rect 239814 285902 239874 285910
rect 239814 285842 240212 285902
rect 188286 285834 188292 285836
rect 84150 285774 188292 285834
rect 78806 285636 78812 285700
rect 78876 285698 78882 285700
rect 79961 285698 80027 285701
rect 78876 285696 80027 285698
rect 78876 285640 79966 285696
rect 80022 285640 80027 285696
rect 78876 285638 80027 285640
rect 78876 285636 78882 285638
rect 79961 285635 80027 285638
rect 81014 285636 81020 285700
rect 81084 285698 81090 285700
rect 81341 285698 81407 285701
rect 81084 285696 81407 285698
rect 81084 285640 81346 285696
rect 81402 285640 81407 285696
rect 81084 285638 81407 285640
rect 81084 285636 81090 285638
rect 81341 285635 81407 285638
rect 83406 285636 83412 285700
rect 83476 285698 83482 285700
rect 84150 285698 84210 285774
rect 188286 285772 188292 285774
rect 188356 285772 188362 285836
rect 83476 285638 84210 285698
rect 83476 285636 83482 285638
rect 86166 285636 86172 285700
rect 86236 285698 86242 285700
rect 86861 285698 86927 285701
rect 86236 285696 86927 285698
rect 86236 285640 86866 285696
rect 86922 285640 86927 285696
rect 86236 285638 86927 285640
rect 86236 285636 86242 285638
rect 86861 285635 86927 285638
rect 88558 285636 88564 285700
rect 88628 285698 88634 285700
rect 89621 285698 89687 285701
rect 88628 285696 89687 285698
rect 88628 285640 89626 285696
rect 89682 285640 89687 285696
rect 88628 285638 89687 285640
rect 88628 285636 88634 285638
rect 89621 285635 89687 285638
rect 93526 285636 93532 285700
rect 93596 285698 93602 285700
rect 93669 285698 93735 285701
rect 93596 285696 93735 285698
rect 93596 285640 93674 285696
rect 93730 285640 93735 285696
rect 93596 285638 93735 285640
rect 93596 285636 93602 285638
rect 93669 285635 93735 285638
rect 101254 285636 101260 285700
rect 101324 285698 101330 285700
rect 102041 285698 102107 285701
rect 101324 285696 102107 285698
rect 101324 285640 102046 285696
rect 102102 285640 102107 285696
rect 101324 285638 102107 285640
rect 101324 285636 101330 285638
rect 102041 285635 102107 285638
rect 103830 285636 103836 285700
rect 103900 285698 103906 285700
rect 104801 285698 104867 285701
rect 106181 285700 106247 285701
rect 106181 285698 106228 285700
rect 103900 285696 104867 285698
rect 103900 285640 104806 285696
rect 104862 285640 104867 285696
rect 103900 285638 104867 285640
rect 106136 285696 106228 285698
rect 106136 285640 106186 285696
rect 106136 285638 106228 285640
rect 103900 285636 103906 285638
rect 104801 285635 104867 285638
rect 106181 285636 106228 285638
rect 106292 285636 106298 285700
rect 120758 285636 120764 285700
rect 120828 285698 120834 285700
rect 121361 285698 121427 285701
rect 120828 285696 121427 285698
rect 120828 285640 121366 285696
rect 121422 285640 121427 285696
rect 120828 285638 121427 285640
rect 120828 285636 120834 285638
rect 106181 285635 106247 285636
rect 121361 285635 121427 285638
rect 138422 285636 138428 285700
rect 138492 285698 138498 285700
rect 139301 285698 139367 285701
rect 138492 285696 139367 285698
rect 138492 285640 139306 285696
rect 139362 285640 139367 285696
rect 138492 285638 139367 285640
rect 138492 285636 138498 285638
rect 139301 285635 139367 285638
rect 140998 285636 141004 285700
rect 141068 285698 141074 285700
rect 142061 285698 142127 285701
rect 141068 285696 142127 285698
rect 141068 285640 142066 285696
rect 142122 285640 142127 285696
rect 141068 285638 142127 285640
rect 141068 285636 141074 285638
rect 142061 285635 142127 285638
rect 143574 285636 143580 285700
rect 143644 285698 143650 285700
rect 144821 285698 144887 285701
rect 143644 285696 144887 285698
rect 143644 285640 144826 285696
rect 144882 285640 144887 285696
rect 143644 285638 144887 285640
rect 143644 285636 143650 285638
rect 144821 285635 144887 285638
rect 145598 285636 145604 285700
rect 145668 285698 145674 285700
rect 146201 285698 146267 285701
rect 145668 285696 146267 285698
rect 145668 285640 146206 285696
rect 146262 285640 146267 285696
rect 145668 285638 146267 285640
rect 145668 285636 145674 285638
rect 146201 285635 146267 285638
rect 148542 285636 148548 285700
rect 148612 285698 148618 285700
rect 148961 285698 149027 285701
rect 148612 285696 149027 285698
rect 148612 285640 148966 285696
rect 149022 285640 149027 285696
rect 148612 285638 149027 285640
rect 148612 285636 148618 285638
rect 148961 285635 149027 285638
rect 151118 285636 151124 285700
rect 151188 285698 151194 285700
rect 151721 285698 151787 285701
rect 151188 285696 151787 285698
rect 151188 285640 151726 285696
rect 151782 285640 151787 285696
rect 151188 285638 151787 285640
rect 151188 285636 151194 285638
rect 151721 285635 151787 285638
rect 154062 285636 154068 285700
rect 154132 285698 154138 285700
rect 154481 285698 154547 285701
rect 154132 285696 154547 285698
rect 154132 285640 154486 285696
rect 154542 285640 154547 285696
rect 154132 285638 154547 285640
rect 154132 285636 154138 285638
rect 154481 285635 154547 285638
rect 156086 285636 156092 285700
rect 156156 285698 156162 285700
rect 157241 285698 157307 285701
rect 156156 285696 157307 285698
rect 156156 285640 157246 285696
rect 157302 285640 157307 285696
rect 156156 285638 157307 285640
rect 156156 285636 156162 285638
rect 157241 285635 157307 285638
rect 583520 285276 584960 285516
rect 96153 285156 96219 285157
rect 113817 285156 113883 285157
rect 123569 285156 123635 285157
rect 128721 285156 128787 285157
rect 96102 285092 96108 285156
rect 96172 285154 96219 285156
rect 96172 285152 96264 285154
rect 96214 285096 96264 285152
rect 96172 285094 96264 285096
rect 96172 285092 96219 285094
rect 113766 285092 113772 285156
rect 113836 285154 113883 285156
rect 113836 285152 113928 285154
rect 113878 285096 113928 285152
rect 113836 285094 113928 285096
rect 113836 285092 113883 285094
rect 123518 285092 123524 285156
rect 123588 285154 123635 285156
rect 123588 285152 123680 285154
rect 123630 285096 123680 285152
rect 123588 285094 123680 285096
rect 123588 285092 123635 285094
rect 128670 285092 128676 285156
rect 128740 285154 128787 285156
rect 128740 285152 128832 285154
rect 128782 285096 128832 285152
rect 128740 285094 128832 285096
rect 128740 285092 128787 285094
rect 96153 285091 96219 285092
rect 113817 285091 113883 285092
rect 123569 285091 123635 285092
rect 128721 285091 128787 285092
rect 98545 285020 98611 285021
rect 118601 285020 118667 285021
rect 98494 284956 98500 285020
rect 98564 285018 98611 285020
rect 98564 285016 98656 285018
rect 98606 284960 98656 285016
rect 98564 284958 98656 284960
rect 98564 284956 98611 284958
rect 118550 284956 118556 285020
rect 118620 285018 118667 285020
rect 118620 285016 118712 285018
rect 118662 284960 118712 285016
rect 118620 284958 118712 284960
rect 118620 284956 118667 284958
rect 98545 284955 98611 284956
rect 118601 284955 118667 284956
rect 91185 284884 91251 284885
rect 91134 284820 91140 284884
rect 91204 284882 91251 284884
rect 91204 284880 91296 284882
rect 91246 284824 91296 284880
rect 91204 284822 91296 284824
rect 91204 284820 91251 284822
rect 91185 284819 91251 284820
rect 239814 284754 240212 284814
rect 237373 284746 237439 284749
rect 239814 284746 239874 284754
rect 237373 284744 239874 284746
rect 237373 284688 237378 284744
rect 237434 284688 239874 284744
rect 237373 284686 239874 284688
rect 237373 284683 237439 284686
rect 180701 284068 180767 284069
rect 180701 284066 180748 284068
rect 180656 284064 180748 284066
rect 180812 284066 180818 284068
rect 180656 284008 180706 284064
rect 180656 284006 180748 284008
rect 180701 284004 180748 284006
rect 180812 284006 180894 284066
rect 180812 284004 180818 284006
rect 180701 284003 180767 284004
rect 239814 283802 240212 283862
rect 237465 283794 237531 283797
rect 239814 283794 239874 283802
rect 237465 283792 239874 283794
rect 237465 283736 237470 283792
rect 237526 283736 239874 283792
rect 237465 283734 239874 283736
rect 237465 283731 237531 283734
rect 237373 282842 237439 282845
rect 237373 282840 239874 282842
rect 237373 282784 237378 282840
rect 237434 282784 239874 282840
rect 237373 282782 239874 282784
rect 237373 282779 237439 282782
rect 239814 282774 239874 282782
rect 239814 282714 240212 282774
rect 239814 281762 240212 281822
rect 237373 281754 237439 281757
rect 239814 281754 239874 281762
rect 237373 281752 239874 281754
rect 237373 281696 237378 281752
rect 237434 281696 239874 281752
rect 237373 281694 239874 281696
rect 237373 281691 237439 281694
rect 239814 280674 240212 280734
rect 237465 280666 237531 280669
rect 239814 280666 239874 280674
rect 237465 280664 239874 280666
rect 237465 280608 237470 280664
rect 237526 280608 239874 280664
rect 237465 280606 239874 280608
rect 237465 280603 237531 280606
rect -960 279972 480 280212
rect 237373 279850 237439 279853
rect 237373 279848 239874 279850
rect 237373 279792 237378 279848
rect 237434 279792 239874 279848
rect 237373 279790 239874 279792
rect 237373 279787 237439 279790
rect 239814 279782 239874 279790
rect 239814 279722 240212 279782
rect 186588 279170 187250 279220
rect 189073 279170 189139 279173
rect 186588 279168 189139 279170
rect 186588 279160 189078 279168
rect 187190 279112 189078 279160
rect 189134 279112 189139 279168
rect 187190 279110 189139 279112
rect 189073 279107 189139 279110
rect 239814 278634 240212 278694
rect 238293 278626 238359 278629
rect 239814 278626 239874 278634
rect 238293 278624 239874 278626
rect 238293 278568 238298 278624
rect 238354 278568 239874 278624
rect 238293 278566 239874 278568
rect 238293 278563 238359 278566
rect 239814 277682 240212 277742
rect 238150 277612 238156 277676
rect 238220 277674 238226 277676
rect 239814 277674 239874 277682
rect 238220 277614 239874 277674
rect 238220 277612 238226 277614
rect 238661 276858 238727 276861
rect 238661 276856 239874 276858
rect 238661 276800 238666 276856
rect 238722 276800 239874 276856
rect 238661 276798 239874 276800
rect 238661 276795 238727 276798
rect 239814 276790 239874 276798
rect 239814 276730 240212 276790
rect 239814 275642 240212 275702
rect 237465 275634 237531 275637
rect 239814 275634 239874 275642
rect 237465 275632 239874 275634
rect 237465 275576 237470 275632
rect 237526 275576 239874 275632
rect 237465 275574 239874 275576
rect 237465 275571 237531 275574
rect 237373 274818 237439 274821
rect 237373 274816 239874 274818
rect 237373 274760 237378 274816
rect 237434 274760 239874 274816
rect 237373 274758 239874 274760
rect 237373 274755 237439 274758
rect 239814 274750 239874 274758
rect 239814 274690 240212 274750
rect 237373 273730 237439 273733
rect 237373 273728 239874 273730
rect 237373 273672 237378 273728
rect 237434 273672 239874 273728
rect 237373 273670 239874 273672
rect 237373 273667 237439 273670
rect 239814 273662 239874 273670
rect 239814 273602 240212 273662
rect 239814 272650 240212 272710
rect 237373 272642 237439 272645
rect 239814 272642 239874 272650
rect 237373 272640 239874 272642
rect 237373 272584 237378 272640
rect 237434 272584 239874 272640
rect 237373 272582 239874 272584
rect 237373 272579 237439 272582
rect 580165 272234 580231 272237
rect 583520 272234 584960 272324
rect 580165 272232 584960 272234
rect 580165 272176 580170 272232
rect 580226 272176 584960 272232
rect 580165 272174 584960 272176
rect 580165 272171 580231 272174
rect 583520 272084 584960 272174
rect 239814 271562 240212 271622
rect 239814 271282 239874 271562
rect 219390 271222 239874 271282
rect 186814 270540 186820 270604
rect 186884 270602 186890 270604
rect 219390 270602 219450 271222
rect 238109 270738 238175 270741
rect 238109 270736 239874 270738
rect 238109 270680 238114 270736
rect 238170 270680 239874 270736
rect 238109 270678 239874 270680
rect 238109 270675 238175 270678
rect 239814 270670 239874 270678
rect 239814 270610 240212 270670
rect 186884 270542 219450 270602
rect 186884 270540 186890 270542
rect 239814 269522 240212 269582
rect 237373 269514 237439 269517
rect 239814 269514 239874 269522
rect 237373 269512 239874 269514
rect 237373 269456 237378 269512
rect 237434 269456 239874 269512
rect 237373 269454 239874 269456
rect 237373 269451 237439 269454
rect 239814 268570 240212 268630
rect 238334 268500 238340 268564
rect 238404 268562 238410 268564
rect 239814 268562 239874 268570
rect 238404 268502 239874 268562
rect 238404 268500 238410 268502
rect 238569 267610 238635 267613
rect 238569 267608 239874 267610
rect 238569 267552 238574 267608
rect 238630 267552 239874 267608
rect 238569 267550 239874 267552
rect 238569 267547 238635 267550
rect 239814 267542 239874 267550
rect 239814 267482 240212 267542
rect -960 267052 480 267292
rect 239814 266530 240212 266590
rect 238109 266522 238175 266525
rect 239814 266522 239874 266530
rect 238109 266520 239874 266522
rect 238109 266464 238114 266520
rect 238170 266464 239874 266520
rect 238109 266462 239874 266464
rect 238109 266459 238175 266462
rect 239814 265578 240212 265638
rect 237373 265570 237439 265573
rect 239814 265570 239874 265578
rect 237373 265568 239874 265570
rect 237373 265512 237378 265568
rect 237434 265512 239874 265568
rect 237373 265510 239874 265512
rect 237373 265507 237439 265510
rect 238385 264618 238451 264621
rect 238385 264616 239874 264618
rect 238385 264560 238390 264616
rect 238446 264560 239874 264616
rect 238385 264558 239874 264560
rect 238385 264555 238451 264558
rect 239814 264550 239874 264558
rect 239814 264490 240212 264550
rect 239814 263538 240212 263598
rect 237373 263530 237439 263533
rect 239814 263530 239874 263538
rect 237373 263528 239874 263530
rect 237373 263472 237378 263528
rect 237434 263472 239874 263528
rect 237373 263470 239874 263472
rect 237373 263467 237439 263470
rect 239814 262450 240212 262510
rect 238518 262380 238524 262444
rect 238588 262442 238594 262444
rect 239814 262442 239874 262450
rect 238588 262382 239874 262442
rect 238588 262380 238594 262382
rect 238201 261626 238267 261629
rect 238201 261624 239874 261626
rect 238201 261568 238206 261624
rect 238262 261568 239874 261624
rect 238201 261566 239874 261568
rect 238201 261563 238267 261566
rect 239814 261558 239874 261566
rect 239814 261498 240212 261558
rect 239814 260410 240212 260470
rect 237465 260402 237531 260405
rect 239814 260402 239874 260410
rect 237465 260400 239874 260402
rect 237465 260344 237470 260400
rect 237526 260344 239874 260400
rect 237465 260342 239874 260344
rect 237465 260339 237531 260342
rect 237373 259586 237439 259589
rect 237373 259584 239874 259586
rect 237373 259528 237378 259584
rect 237434 259528 239874 259584
rect 237373 259526 239874 259528
rect 237373 259523 237439 259526
rect 239814 259518 239874 259526
rect 239814 259458 240212 259518
rect 580901 258906 580967 258909
rect 583520 258906 584960 258996
rect 580901 258904 584960 258906
rect 580901 258848 580906 258904
rect 580962 258848 584960 258904
rect 580901 258846 584960 258848
rect 580901 258843 580967 258846
rect 583520 258756 584960 258846
rect 237373 258498 237439 258501
rect 237373 258496 239874 258498
rect 237373 258440 237378 258496
rect 237434 258440 239874 258496
rect 237373 258438 239874 258440
rect 237373 258435 237439 258438
rect 239814 258430 239874 258438
rect 239814 258370 240212 258430
rect 239814 257418 240212 257478
rect 238201 257410 238267 257413
rect 239814 257410 239874 257418
rect 238201 257408 239874 257410
rect 238201 257352 238206 257408
rect 238262 257352 239874 257408
rect 238201 257350 239874 257352
rect 238201 257347 238267 257350
rect 239814 256330 240212 256390
rect 237373 256322 237439 256325
rect 239814 256322 239874 256330
rect 237373 256320 239874 256322
rect 237373 256264 237378 256320
rect 237434 256264 239874 256320
rect 237373 256262 239874 256264
rect 237373 256259 237439 256262
rect 237465 255506 237531 255509
rect 237465 255504 239874 255506
rect 237465 255448 237470 255504
rect 237526 255448 239874 255504
rect 237465 255446 239874 255448
rect 237465 255443 237531 255446
rect 239814 255438 239874 255446
rect 239814 255378 240212 255438
rect 239814 254426 240212 254486
rect 237373 254418 237439 254421
rect 239814 254418 239874 254426
rect 237373 254416 239874 254418
rect 237373 254360 237378 254416
rect 237434 254360 239874 254416
rect 237373 254358 239874 254360
rect 237373 254355 237439 254358
rect -960 254146 480 254236
rect 3969 254146 4035 254149
rect -960 254144 4035 254146
rect -960 254088 3974 254144
rect 4030 254088 4035 254144
rect -960 254086 4035 254088
rect -960 253996 480 254086
rect 3969 254083 4035 254086
rect 239814 253338 240212 253398
rect 237465 253330 237531 253333
rect 239814 253330 239874 253338
rect 237465 253328 239874 253330
rect 237465 253272 237470 253328
rect 237526 253272 239874 253328
rect 237465 253270 239874 253272
rect 237465 253267 237531 253270
rect 237373 252514 237439 252517
rect 237373 252512 239874 252514
rect 237373 252456 237378 252512
rect 237434 252456 239874 252512
rect 237373 252454 239874 252456
rect 237373 252451 237439 252454
rect 239814 252446 239874 252454
rect 239814 252386 240212 252446
rect 239814 251298 240212 251358
rect 238385 251290 238451 251293
rect 239814 251290 239874 251298
rect 238385 251288 239874 251290
rect 238385 251232 238390 251288
rect 238446 251232 239874 251288
rect 238385 251230 239874 251232
rect 238385 251227 238451 251230
rect 239814 250346 240212 250406
rect 237373 250338 237439 250341
rect 239814 250338 239874 250346
rect 237373 250336 239874 250338
rect 237373 250280 237378 250336
rect 237434 250280 239874 250336
rect 237373 250278 239874 250280
rect 237373 250275 237439 250278
rect 237373 247346 237439 247349
rect 237373 247344 239874 247346
rect 237373 247288 237378 247344
rect 237434 247288 239874 247344
rect 237373 247286 239874 247288
rect 237373 247283 237439 247286
rect 239814 247278 239874 247286
rect 239814 247218 240212 247278
rect 239814 246266 240212 246326
rect 237373 246258 237439 246261
rect 239814 246258 239874 246266
rect 237373 246256 239874 246258
rect 237373 246200 237378 246256
rect 237434 246200 239874 246256
rect 237373 246198 239874 246200
rect 237373 246195 237439 246198
rect 583520 245428 584960 245668
rect 239814 245178 240212 245238
rect 237373 245170 237439 245173
rect 239814 245170 239874 245178
rect 237373 245168 239874 245170
rect 237373 245112 237378 245168
rect 237434 245112 239874 245168
rect 237373 245110 239874 245112
rect 237373 245107 237439 245110
rect 237373 242314 237439 242317
rect 237373 242312 239874 242314
rect 237373 242256 237378 242312
rect 237434 242256 239874 242312
rect 237373 242254 239874 242256
rect 237373 242251 237439 242254
rect 239814 242246 239874 242254
rect 239814 242186 240212 242246
rect 239814 241234 240212 241294
rect 238569 241226 238635 241229
rect 239814 241226 239874 241234
rect 238569 241224 239874 241226
rect -960 241090 480 241180
rect 238569 241168 238574 241224
rect 238630 241168 239874 241224
rect 238569 241166 239874 241168
rect 238569 241163 238635 241166
rect 3233 241090 3299 241093
rect -960 241088 3299 241090
rect -960 241032 3238 241088
rect 3294 241032 3299 241088
rect -960 241030 3299 241032
rect -960 240940 480 241030
rect 3233 241027 3299 241030
rect 237373 240274 237439 240277
rect 237373 240272 239874 240274
rect 237373 240216 237378 240272
rect 237434 240216 239874 240272
rect 237373 240214 239874 240216
rect 237373 240211 237439 240214
rect 239814 240206 239874 240214
rect 239814 240146 240212 240206
rect 237373 237282 237439 237285
rect 237373 237280 239874 237282
rect 237373 237224 237378 237280
rect 237434 237224 239874 237280
rect 237373 237222 239874 237224
rect 237373 237219 237439 237222
rect 239814 237214 239874 237222
rect 239814 237154 240212 237214
rect 48129 236874 48195 236877
rect 49374 236874 50048 236924
rect 48129 236872 50048 236874
rect 48129 236816 48134 236872
rect 48190 236864 50048 236872
rect 48190 236816 49434 236864
rect 48129 236814 49434 236816
rect 48129 236811 48195 236814
rect 239814 236066 240212 236126
rect 237373 236058 237439 236061
rect 239814 236058 239874 236066
rect 237373 236056 239874 236058
rect 237373 236000 237378 236056
rect 237434 236000 239874 236056
rect 237373 235998 239874 236000
rect 237373 235995 237439 235998
rect 47945 235922 48011 235925
rect 49374 235922 50048 235972
rect 47945 235920 50048 235922
rect 47945 235864 47950 235920
rect 48006 235912 50048 235920
rect 48006 235864 49434 235912
rect 47945 235862 49434 235864
rect 47945 235859 48011 235862
rect 239814 235114 240212 235174
rect 186998 234636 187004 234700
rect 187068 234698 187074 234700
rect 239814 234698 239874 235114
rect 187068 234638 239874 234698
rect 187068 234636 187074 234638
rect 48037 233746 48103 233749
rect 49374 233746 50048 233796
rect 48037 233744 50048 233746
rect 48037 233688 48042 233744
rect 48098 233736 50048 233744
rect 48098 233688 49434 233736
rect 48037 233686 49434 233688
rect 48037 233683 48103 233686
rect 47761 232794 47827 232797
rect 49374 232794 50048 232844
rect 47761 232792 50048 232794
rect 47761 232736 47766 232792
rect 47822 232784 50048 232792
rect 47822 232736 49434 232784
rect 47761 232734 49434 232736
rect 47761 232731 47827 232734
rect 580165 232386 580231 232389
rect 583520 232386 584960 232476
rect 580165 232384 584960 232386
rect 580165 232328 580170 232384
rect 580226 232328 584960 232384
rect 580165 232326 584960 232328
rect 580165 232323 580231 232326
rect 238477 232250 238543 232253
rect 238477 232248 239874 232250
rect 238477 232192 238482 232248
rect 238538 232192 239874 232248
rect 583520 232236 584960 232326
rect 238477 232190 239874 232192
rect 238477 232187 238543 232190
rect 239814 232182 239874 232190
rect 239814 232122 240212 232182
rect 47669 231026 47735 231029
rect 49374 231026 50048 231076
rect 239814 231034 240212 231094
rect 47669 231024 50048 231026
rect 47669 230968 47674 231024
rect 47730 231016 50048 231024
rect 237373 231026 237439 231029
rect 239814 231026 239874 231034
rect 237373 231024 239874 231026
rect 47730 230968 49434 231016
rect 47669 230966 49434 230968
rect 237373 230968 237378 231024
rect 237434 230968 239874 231024
rect 237373 230966 239874 230968
rect 47669 230963 47735 230966
rect 237373 230963 237439 230966
rect 239814 230082 240212 230142
rect 238477 230074 238543 230077
rect 239814 230074 239874 230082
rect 238477 230072 239874 230074
rect 238477 230016 238482 230072
rect 238538 230016 239874 230072
rect 238477 230014 239874 230016
rect 238477 230011 238543 230014
rect 47853 229938 47919 229941
rect 49374 229938 50048 229988
rect 47853 229936 50048 229938
rect 47853 229880 47858 229936
rect 47914 229928 50048 229936
rect 47914 229880 49434 229928
rect 47853 229878 49434 229880
rect 47853 229875 47919 229878
rect 239814 228994 240212 229054
rect 237465 228986 237531 228989
rect 239814 228986 239874 228994
rect 237465 228984 239874 228986
rect 237465 228928 237470 228984
rect 237526 228928 239874 228984
rect 237465 228926 239874 228928
rect 237465 228923 237531 228926
rect 49509 228220 49575 228223
rect 49509 228218 50048 228220
rect 49509 228162 49514 228218
rect 49570 228162 50048 228218
rect 49509 228160 50048 228162
rect 49509 228157 49575 228160
rect -960 227884 480 228124
rect 239814 228042 240212 228102
rect 237373 228034 237439 228037
rect 239814 228034 239874 228042
rect 237373 228032 239874 228034
rect 237373 227976 237378 228032
rect 237434 227976 239874 228032
rect 237373 227974 239874 227976
rect 237373 227971 237439 227974
rect 237373 227082 237439 227085
rect 237373 227080 239874 227082
rect 237373 227024 237378 227080
rect 237434 227024 239874 227080
rect 237373 227022 239874 227024
rect 237373 227019 237439 227022
rect 239814 227014 239874 227022
rect 239814 226954 240212 227014
rect 239814 226002 240212 226062
rect 237373 225994 237439 225997
rect 239814 225994 239874 226002
rect 237373 225992 239874 225994
rect 237373 225936 237378 225992
rect 237434 225936 239874 225992
rect 237373 225934 239874 225936
rect 237373 225931 237439 225934
rect 238661 225042 238727 225045
rect 238661 225040 239874 225042
rect 238661 224984 238666 225040
rect 238722 224984 239874 225040
rect 238661 224982 239874 224984
rect 238661 224979 238727 224982
rect 239814 224970 239874 224982
rect 239814 224910 240242 224970
rect 239814 223962 240212 224022
rect 237373 223954 237439 223957
rect 239814 223954 239874 223962
rect 237373 223952 239874 223954
rect 237373 223896 237378 223952
rect 237434 223896 239874 223952
rect 237373 223894 239874 223896
rect 237373 223891 237439 223894
rect 239814 223010 240212 223070
rect 237925 223002 237991 223005
rect 239814 223002 239874 223010
rect 237925 223000 239874 223002
rect 237925 222944 237930 223000
rect 237986 222944 239874 223000
rect 237925 222942 239874 222944
rect 237925 222939 237991 222942
rect 188470 222804 188476 222868
rect 188540 222866 188546 222868
rect 238293 222866 238359 222869
rect 188540 222864 238359 222866
rect 188540 222808 238298 222864
rect 238354 222808 238359 222864
rect 188540 222806 238359 222808
rect 188540 222804 188546 222806
rect 238293 222803 238359 222806
rect 237373 222050 237439 222053
rect 237373 222048 239874 222050
rect 237373 221992 237378 222048
rect 237434 221992 239874 222048
rect 237373 221990 239874 221992
rect 237373 221987 237439 221990
rect 239814 221982 239874 221990
rect 239814 221922 240212 221982
rect 239814 220970 240212 221030
rect 237373 220962 237439 220965
rect 239814 220962 239874 220970
rect 237373 220960 239874 220962
rect 237373 220904 237378 220960
rect 237434 220904 239874 220960
rect 237373 220902 239874 220904
rect 237373 220899 237439 220902
rect 239814 219882 240212 219942
rect 238293 219874 238359 219877
rect 239814 219874 239874 219882
rect 238293 219872 239874 219874
rect 238293 219816 238298 219872
rect 238354 219816 239874 219872
rect 238293 219814 239874 219816
rect 238293 219811 238359 219814
rect 186588 219330 187250 219380
rect 189073 219330 189139 219333
rect 186588 219328 189139 219330
rect 186588 219320 189078 219328
rect 187190 219272 189078 219320
rect 189134 219272 189139 219328
rect 187190 219270 189139 219272
rect 189073 219267 189139 219270
rect 580165 219058 580231 219061
rect 583520 219058 584960 219148
rect 580165 219056 584960 219058
rect 580165 219000 580170 219056
rect 580226 219000 584960 219056
rect 580165 218998 584960 219000
rect 580165 218995 580231 218998
rect 239814 218930 240212 218990
rect 237373 218922 237439 218925
rect 239814 218922 239874 218930
rect 237373 218920 239874 218922
rect 237373 218864 237378 218920
rect 237434 218864 239874 218920
rect 583520 218908 584960 218998
rect 237373 218862 239874 218864
rect 237373 218859 237439 218862
rect 239814 217842 240212 217902
rect 237373 217834 237439 217837
rect 239814 217834 239874 217842
rect 237373 217832 239874 217834
rect 237373 217776 237378 217832
rect 237434 217776 239874 217832
rect 237373 217774 239874 217776
rect 237373 217771 237439 217774
rect 186588 217698 187250 217748
rect 189073 217698 189139 217701
rect 186588 217696 189139 217698
rect 186588 217688 189078 217696
rect 187190 217640 189078 217688
rect 189134 217640 189139 217696
rect 187190 217638 189139 217640
rect 189073 217635 189139 217638
rect 238017 217018 238083 217021
rect 238017 217016 239874 217018
rect 238017 216960 238022 217016
rect 238078 216960 239874 217016
rect 238017 216958 239874 216960
rect 238017 216955 238083 216958
rect 239814 216950 239874 216958
rect 239814 216890 240212 216950
rect 186588 216338 187250 216388
rect 189165 216338 189231 216341
rect 186588 216336 189231 216338
rect 186588 216328 189170 216336
rect 187190 216280 189170 216328
rect 189226 216280 189231 216336
rect 187190 216278 189231 216280
rect 189165 216275 189231 216278
rect 239814 215802 240212 215862
rect 237373 215794 237439 215797
rect 239814 215794 239874 215802
rect 237373 215792 239874 215794
rect 237373 215736 237378 215792
rect 237434 215736 239874 215792
rect 237373 215734 239874 215736
rect 237373 215731 237439 215734
rect -960 214828 480 215068
rect 186588 214842 187250 214892
rect 239814 214850 240212 214910
rect 190453 214842 190519 214845
rect 186588 214840 190519 214842
rect 186588 214832 190458 214840
rect 187190 214784 190458 214832
rect 190514 214784 190519 214840
rect 187190 214782 190519 214784
rect 190453 214779 190519 214782
rect 237465 214842 237531 214845
rect 239814 214842 239874 214850
rect 237465 214840 239874 214842
rect 237465 214784 237470 214840
rect 237526 214784 239874 214840
rect 237465 214782 239874 214784
rect 237465 214779 237531 214782
rect 237373 213890 237439 213893
rect 237373 213888 239874 213890
rect 237373 213832 237378 213888
rect 237434 213832 239874 213888
rect 237373 213830 239874 213832
rect 237373 213827 237439 213830
rect 239814 213822 239874 213830
rect 239814 213762 240212 213822
rect 189073 213754 189139 213757
rect 187190 213752 189139 213754
rect 187190 213696 189078 213752
rect 189134 213696 189139 213752
rect 187190 213694 189139 213696
rect 187190 213668 187250 213694
rect 189073 213691 189139 213694
rect 186588 213608 187250 213668
rect 239814 212810 240212 212870
rect 237373 212802 237439 212805
rect 239814 212802 239874 212810
rect 237373 212800 239874 212802
rect 237373 212744 237378 212800
rect 237434 212744 239874 212800
rect 237373 212742 239874 212744
rect 237373 212739 237439 212742
rect 237465 211986 237531 211989
rect 237465 211984 239874 211986
rect 237465 211928 237470 211984
rect 237526 211928 239874 211984
rect 237465 211926 239874 211928
rect 237465 211923 237531 211926
rect 239814 211918 239874 211926
rect 239814 211858 240212 211918
rect 239814 210770 240212 210830
rect 237465 210762 237531 210765
rect 239814 210762 239874 210770
rect 237465 210760 239874 210762
rect 237465 210704 237470 210760
rect 237526 210704 239874 210760
rect 237465 210702 239874 210704
rect 237465 210699 237531 210702
rect 49325 209946 49391 209949
rect 49742 209946 50048 209996
rect 49325 209944 50048 209946
rect 49325 209888 49330 209944
rect 49386 209936 50048 209944
rect 49386 209888 49802 209936
rect 49325 209886 49802 209888
rect 49325 209883 49391 209886
rect 239814 209818 240212 209878
rect 237373 209810 237439 209813
rect 239814 209810 239874 209818
rect 237373 209808 239874 209810
rect 237373 209752 237378 209808
rect 237434 209752 239874 209808
rect 237373 209750 239874 209752
rect 237373 209747 237439 209750
rect 237465 208858 237531 208861
rect 237465 208856 239874 208858
rect 237465 208800 237470 208856
rect 237526 208800 239874 208856
rect 237465 208798 239874 208800
rect 237465 208795 237531 208798
rect 239814 208790 239874 208798
rect 239814 208730 240212 208790
rect 49601 208364 49667 208367
rect 49601 208362 50048 208364
rect 49601 208306 49606 208362
rect 49662 208306 50048 208362
rect 49601 208304 50048 208306
rect 49601 208301 49667 208304
rect 49417 208092 49483 208095
rect 49417 208090 50048 208092
rect 49417 208034 49422 208090
rect 49478 208034 50048 208090
rect 49417 208032 50048 208034
rect 49417 208029 49483 208032
rect 239814 207778 240212 207838
rect 237373 207770 237439 207773
rect 239814 207770 239874 207778
rect 237373 207768 239874 207770
rect 237373 207712 237378 207768
rect 237434 207712 239874 207768
rect 237373 207710 239874 207712
rect 237373 207707 237439 207710
rect 239814 206690 240212 206750
rect 237373 206682 237439 206685
rect 239814 206682 239874 206690
rect 237373 206680 239874 206682
rect 237373 206624 237378 206680
rect 237434 206624 239874 206680
rect 237373 206622 239874 206624
rect 237373 206619 237439 206622
rect 237465 205866 237531 205869
rect 237465 205864 239874 205866
rect 237465 205808 237470 205864
rect 237526 205808 239874 205864
rect 237465 205806 239874 205808
rect 237465 205803 237531 205806
rect 239814 205798 239874 205806
rect 239814 205738 240212 205798
rect 583520 205580 584960 205820
rect 239814 204650 240212 204710
rect 238017 204642 238083 204645
rect 239814 204642 239874 204650
rect 238017 204640 239874 204642
rect 238017 204584 238022 204640
rect 238078 204584 239874 204640
rect 238017 204582 239874 204584
rect 238017 204579 238083 204582
rect 239814 203698 240212 203758
rect 237833 203690 237899 203693
rect 239814 203690 239874 203698
rect 237833 203688 239874 203690
rect 237833 203632 237838 203688
rect 237894 203632 239874 203688
rect 237833 203630 239874 203632
rect 237833 203627 237899 203630
rect 237373 202738 237439 202741
rect 237373 202736 239874 202738
rect 237373 202680 237378 202736
rect 237434 202680 239874 202736
rect 237373 202678 239874 202680
rect 237373 202675 237439 202678
rect 239814 202670 239874 202678
rect 239814 202610 240212 202670
rect -960 201922 480 202012
rect 4061 201922 4127 201925
rect -960 201920 4127 201922
rect -960 201864 4066 201920
rect 4122 201864 4127 201920
rect -960 201862 4127 201864
rect -960 201772 480 201862
rect 4061 201859 4127 201862
rect 239814 201658 240212 201718
rect 237373 201650 237439 201653
rect 239814 201650 239874 201658
rect 237373 201648 239874 201650
rect 237373 201592 237378 201648
rect 237434 201592 239874 201648
rect 237373 201590 239874 201592
rect 237373 201587 237439 201590
rect 238334 200834 238340 200836
rect 219390 200774 238340 200834
rect 187550 200636 187556 200700
rect 187620 200698 187626 200700
rect 219390 200698 219450 200774
rect 238334 200772 238340 200774
rect 238404 200772 238410 200836
rect 239814 200706 240212 200766
rect 187620 200638 219450 200698
rect 237373 200698 237439 200701
rect 239814 200698 239874 200706
rect 237373 200696 239874 200698
rect 237373 200640 237378 200696
rect 237434 200640 239874 200696
rect 237373 200638 239874 200640
rect 187620 200636 187626 200638
rect 237373 200635 237439 200638
rect 48129 199882 48195 199885
rect 235809 199882 235875 199885
rect 48129 199880 235875 199882
rect 48129 199824 48134 199880
rect 48190 199824 235814 199880
rect 235870 199824 235875 199880
rect 48129 199822 235875 199824
rect 48129 199819 48195 199822
rect 235809 199819 235875 199822
rect 47761 199746 47827 199749
rect 190361 199746 190427 199749
rect 47761 199744 190427 199746
rect 47761 199688 47766 199744
rect 47822 199688 190366 199744
rect 190422 199688 190427 199744
rect 47761 199686 190427 199688
rect 47761 199683 47827 199686
rect 190361 199683 190427 199686
rect 239814 199618 240212 199678
rect 47669 199610 47735 199613
rect 189625 199610 189691 199613
rect 47669 199608 189691 199610
rect 47669 199552 47674 199608
rect 47730 199552 189630 199608
rect 189686 199552 189691 199608
rect 47669 199550 189691 199552
rect 47669 199547 47735 199550
rect 189625 199547 189691 199550
rect 70577 199476 70643 199477
rect 77753 199476 77819 199477
rect 78857 199476 78923 199477
rect 88609 199476 88675 199477
rect 91185 199476 91251 199477
rect 103697 199476 103763 199477
rect 111057 199476 111123 199477
rect 70526 199474 70532 199476
rect 70486 199414 70532 199474
rect 70596 199472 70643 199476
rect 77702 199474 77708 199476
rect 70638 199416 70643 199472
rect 70526 199412 70532 199414
rect 70596 199412 70643 199416
rect 77662 199414 77708 199474
rect 77772 199472 77819 199476
rect 78806 199474 78812 199476
rect 77814 199416 77819 199472
rect 77702 199412 77708 199414
rect 77772 199412 77819 199416
rect 78766 199414 78812 199474
rect 78876 199472 78923 199476
rect 88558 199474 88564 199476
rect 78918 199416 78923 199472
rect 78806 199412 78812 199414
rect 78876 199412 78923 199416
rect 88518 199414 88564 199474
rect 88628 199472 88675 199476
rect 91134 199474 91140 199476
rect 88670 199416 88675 199472
rect 88558 199412 88564 199414
rect 88628 199412 88675 199416
rect 91094 199414 91140 199474
rect 91204 199472 91251 199476
rect 103646 199474 103652 199476
rect 91246 199416 91251 199472
rect 91134 199412 91140 199414
rect 91204 199412 91251 199416
rect 103606 199414 103652 199474
rect 103716 199472 103763 199476
rect 111006 199474 111012 199476
rect 103758 199416 103763 199472
rect 103646 199412 103652 199414
rect 103716 199412 103763 199416
rect 110966 199414 111012 199474
rect 111076 199472 111123 199476
rect 111118 199416 111123 199472
rect 111006 199412 111012 199414
rect 111076 199412 111123 199416
rect 70577 199411 70643 199412
rect 77753 199411 77819 199412
rect 78857 199411 78923 199412
rect 88609 199411 88675 199412
rect 91185 199411 91251 199412
rect 103697 199411 103763 199412
rect 111057 199411 111123 199412
rect 188286 199140 188292 199204
rect 188356 199202 188362 199204
rect 239814 199202 239874 199618
rect 188356 199142 239874 199202
rect 188356 199140 188362 199142
rect 98678 199004 98684 199068
rect 98748 199066 98754 199068
rect 191189 199066 191255 199069
rect 98748 199064 191255 199066
rect 98748 199008 191194 199064
rect 191250 199008 191255 199064
rect 98748 199006 191255 199008
rect 98748 199004 98754 199006
rect 191189 199003 191255 199006
rect 96470 198868 96476 198932
rect 96540 198930 96546 198932
rect 189809 198930 189875 198933
rect 96540 198928 189875 198930
rect 96540 198872 189814 198928
rect 189870 198872 189875 198928
rect 96540 198870 189875 198872
rect 96540 198868 96546 198870
rect 189809 198867 189875 198870
rect 136030 198732 136036 198796
rect 136100 198794 136106 198796
rect 232865 198794 232931 198797
rect 136100 198792 232931 198794
rect 136100 198736 232870 198792
rect 232926 198736 232931 198792
rect 136100 198734 232931 198736
rect 136100 198732 136106 198734
rect 232865 198731 232931 198734
rect 239998 198726 240242 198760
rect 239814 198700 240242 198726
rect 239814 198666 240058 198700
rect 240182 198696 240242 198700
rect 71865 198660 71931 198661
rect 75545 198660 75611 198661
rect 71814 198658 71820 198660
rect 71774 198598 71820 198658
rect 71884 198656 71931 198660
rect 75494 198658 75500 198660
rect 71926 198600 71931 198656
rect 71814 198596 71820 198598
rect 71884 198596 71931 198600
rect 75454 198598 75500 198658
rect 75564 198656 75611 198660
rect 75606 198600 75611 198656
rect 75494 198596 75500 198598
rect 75564 198596 75611 198600
rect 76598 198596 76604 198660
rect 76668 198658 76674 198660
rect 76833 198658 76899 198661
rect 80145 198660 80211 198661
rect 80094 198658 80100 198660
rect 76668 198656 76899 198658
rect 76668 198600 76838 198656
rect 76894 198600 76899 198656
rect 76668 198598 76899 198600
rect 80054 198598 80100 198658
rect 80164 198656 80211 198660
rect 80206 198600 80211 198656
rect 76668 198596 76674 198598
rect 71865 198595 71931 198596
rect 75545 198595 75611 198596
rect 76833 198595 76899 198598
rect 80094 198596 80100 198598
rect 80164 198596 80211 198600
rect 80145 198595 80211 198596
rect 81341 198660 81407 198661
rect 82537 198660 82603 198661
rect 84561 198660 84627 198661
rect 86217 198660 86283 198661
rect 81341 198656 81388 198660
rect 81452 198658 81458 198660
rect 82486 198658 82492 198660
rect 81341 198600 81346 198656
rect 81341 198596 81388 198600
rect 81452 198598 81498 198658
rect 82446 198598 82492 198658
rect 82556 198656 82603 198660
rect 84510 198658 84516 198660
rect 82598 198600 82603 198656
rect 81452 198596 81458 198598
rect 82486 198596 82492 198598
rect 82556 198596 82603 198600
rect 84470 198598 84516 198658
rect 84580 198656 84627 198660
rect 86166 198658 86172 198660
rect 84622 198600 84627 198656
rect 84510 198596 84516 198598
rect 84580 198596 84627 198600
rect 86126 198598 86172 198658
rect 86236 198656 86283 198660
rect 86278 198600 86283 198656
rect 86166 198596 86172 198598
rect 86236 198596 86283 198600
rect 87086 198596 87092 198660
rect 87156 198658 87162 198660
rect 87965 198658 88031 198661
rect 92841 198660 92907 198661
rect 93577 198660 93643 198661
rect 95969 198660 96035 198661
rect 104433 198660 104499 198661
rect 105905 198660 105971 198661
rect 106089 198660 106155 198661
rect 108481 198660 108547 198661
rect 113633 198660 113699 198661
rect 92790 198658 92796 198660
rect 87156 198656 88031 198658
rect 87156 198600 87970 198656
rect 88026 198600 88031 198656
rect 87156 198598 88031 198600
rect 92750 198598 92796 198658
rect 92860 198656 92907 198660
rect 93526 198658 93532 198660
rect 92902 198600 92907 198656
rect 87156 198596 87162 198598
rect 81341 198595 81407 198596
rect 82537 198595 82603 198596
rect 84561 198595 84627 198596
rect 86217 198595 86283 198596
rect 87965 198595 88031 198598
rect 92790 198596 92796 198598
rect 92860 198596 92907 198600
rect 93486 198598 93532 198658
rect 93596 198656 93643 198660
rect 95918 198658 95924 198660
rect 93638 198600 93643 198656
rect 93526 198596 93532 198598
rect 93596 198596 93643 198600
rect 95878 198598 95924 198658
rect 95988 198656 96035 198660
rect 96030 198600 96035 198656
rect 95918 198596 95924 198598
rect 95988 198596 96035 198600
rect 97574 198596 97580 198660
rect 97644 198658 97650 198660
rect 104382 198658 104388 198660
rect 97644 198598 103530 198658
rect 104342 198598 104388 198658
rect 104452 198656 104499 198660
rect 105854 198658 105860 198660
rect 104494 198600 104499 198656
rect 97644 198596 97650 198598
rect 92841 198595 92907 198596
rect 93577 198595 93643 198596
rect 95969 198595 96035 198596
rect 85849 198524 85915 198525
rect 88241 198524 88307 198525
rect 89529 198524 89595 198525
rect 90817 198524 90883 198525
rect 98361 198524 98427 198525
rect 85798 198522 85804 198524
rect 85758 198462 85804 198522
rect 85868 198520 85915 198524
rect 88190 198522 88196 198524
rect 85910 198464 85915 198520
rect 85798 198460 85804 198462
rect 85868 198460 85915 198464
rect 88150 198462 88196 198522
rect 88260 198520 88307 198524
rect 89478 198522 89484 198524
rect 88302 198464 88307 198520
rect 88190 198460 88196 198462
rect 88260 198460 88307 198464
rect 89438 198462 89484 198522
rect 89548 198520 89595 198524
rect 90766 198522 90772 198524
rect 89590 198464 89595 198520
rect 89478 198460 89484 198462
rect 89548 198460 89595 198464
rect 90726 198462 90772 198522
rect 90836 198520 90883 198524
rect 98310 198522 98316 198524
rect 90878 198464 90883 198520
rect 90766 198460 90772 198462
rect 90836 198460 90883 198464
rect 98270 198462 98316 198522
rect 98380 198520 98427 198524
rect 98422 198464 98427 198520
rect 98310 198460 98316 198462
rect 98380 198460 98427 198464
rect 99782 198460 99788 198524
rect 99852 198522 99858 198524
rect 100017 198522 100083 198525
rect 100937 198524 101003 198525
rect 102225 198524 102291 198525
rect 103329 198524 103395 198525
rect 100886 198522 100892 198524
rect 99852 198520 100083 198522
rect 99852 198464 100022 198520
rect 100078 198464 100083 198520
rect 99852 198462 100083 198464
rect 100846 198462 100892 198522
rect 100956 198520 101003 198524
rect 102174 198522 102180 198524
rect 100998 198464 101003 198520
rect 99852 198460 99858 198462
rect 85849 198459 85915 198460
rect 88241 198459 88307 198460
rect 89529 198459 89595 198460
rect 90817 198459 90883 198460
rect 98361 198459 98427 198460
rect 100017 198459 100083 198462
rect 100886 198460 100892 198462
rect 100956 198460 101003 198464
rect 102134 198462 102180 198522
rect 102244 198520 102291 198524
rect 103278 198522 103284 198524
rect 102286 198464 102291 198520
rect 102174 198460 102180 198462
rect 102244 198460 102291 198464
rect 103238 198462 103284 198522
rect 103348 198520 103395 198524
rect 103390 198464 103395 198520
rect 103278 198460 103284 198462
rect 103348 198460 103395 198464
rect 103470 198522 103530 198598
rect 104382 198596 104388 198598
rect 104452 198596 104499 198600
rect 105814 198598 105860 198658
rect 105924 198656 105971 198660
rect 105966 198600 105971 198656
rect 105854 198596 105860 198598
rect 105924 198596 105971 198600
rect 106038 198596 106044 198660
rect 106108 198658 106155 198660
rect 108430 198658 108436 198660
rect 106108 198656 106200 198658
rect 106150 198600 106200 198656
rect 106108 198598 106200 198600
rect 108390 198598 108436 198658
rect 108500 198656 108547 198660
rect 113582 198658 113588 198660
rect 108542 198600 108547 198656
rect 106108 198596 106155 198598
rect 108430 198596 108436 198598
rect 108500 198596 108547 198600
rect 113542 198598 113588 198658
rect 113652 198656 113699 198660
rect 113694 198600 113699 198656
rect 113582 198596 113588 198598
rect 113652 198596 113699 198600
rect 115974 198596 115980 198660
rect 116044 198658 116050 198660
rect 117037 198658 117103 198661
rect 118417 198660 118483 198661
rect 120993 198660 121059 198661
rect 123569 198660 123635 198661
rect 118366 198658 118372 198660
rect 116044 198656 117103 198658
rect 116044 198600 117042 198656
rect 117098 198600 117103 198656
rect 116044 198598 117103 198600
rect 118326 198598 118372 198658
rect 118436 198656 118483 198660
rect 120942 198658 120948 198660
rect 118478 198600 118483 198656
rect 116044 198596 116050 198598
rect 104433 198595 104499 198596
rect 105905 198595 105971 198596
rect 106089 198595 106155 198596
rect 108481 198595 108547 198596
rect 113633 198595 113699 198596
rect 117037 198595 117103 198598
rect 118366 198596 118372 198598
rect 118436 198596 118483 198600
rect 120902 198598 120948 198658
rect 121012 198656 121059 198660
rect 123518 198658 123524 198660
rect 121054 198600 121059 198656
rect 120942 198596 120948 198598
rect 121012 198596 121059 198600
rect 123478 198598 123524 198658
rect 123588 198656 123635 198660
rect 123630 198600 123635 198656
rect 123518 198596 123524 198598
rect 123588 198596 123635 198600
rect 125910 198596 125916 198660
rect 125980 198658 125986 198660
rect 126605 198658 126671 198661
rect 125980 198656 126671 198658
rect 125980 198600 126610 198656
rect 126666 198600 126671 198656
rect 125980 198598 126671 198600
rect 125980 198596 125986 198598
rect 118417 198595 118483 198596
rect 120993 198595 121059 198596
rect 123569 198595 123635 198596
rect 126605 198595 126671 198598
rect 128486 198596 128492 198660
rect 128556 198658 128562 198660
rect 128905 198658 128971 198661
rect 146017 198660 146083 198661
rect 153377 198660 153443 198661
rect 173433 198660 173499 198661
rect 145966 198658 145972 198660
rect 128556 198656 128971 198658
rect 128556 198600 128910 198656
rect 128966 198600 128971 198656
rect 128556 198598 128971 198600
rect 145926 198598 145972 198658
rect 146036 198656 146083 198660
rect 153326 198658 153332 198660
rect 146078 198600 146083 198656
rect 128556 198596 128562 198598
rect 128905 198595 128971 198598
rect 145966 198596 145972 198598
rect 146036 198596 146083 198600
rect 153286 198598 153332 198658
rect 153396 198656 153443 198660
rect 173382 198658 173388 198660
rect 153438 198600 153443 198656
rect 153326 198596 153332 198598
rect 153396 198596 153443 198600
rect 173342 198598 173388 198658
rect 173452 198656 173499 198660
rect 173494 198600 173499 198656
rect 173382 198596 173388 198598
rect 173452 198596 173499 198600
rect 146017 198595 146083 198596
rect 153377 198595 153443 198596
rect 173433 198595 173499 198596
rect 237465 198658 237531 198661
rect 239814 198658 239874 198666
rect 237465 198656 239874 198658
rect 237465 198600 237470 198656
rect 237526 198600 239874 198656
rect 237465 198598 239874 198600
rect 237465 198595 237531 198598
rect 238150 198522 238156 198524
rect 103470 198462 238156 198522
rect 238150 198460 238156 198462
rect 238220 198460 238226 198524
rect 100937 198459 101003 198460
rect 102225 198459 102291 198460
rect 103329 198459 103395 198460
rect 73102 198324 73108 198388
rect 73172 198386 73178 198388
rect 73429 198386 73495 198389
rect 73172 198384 73495 198386
rect 73172 198328 73434 198384
rect 73490 198328 73495 198384
rect 73172 198326 73495 198328
rect 73172 198324 73178 198326
rect 73429 198323 73495 198326
rect 83406 198324 83412 198388
rect 83476 198386 83482 198388
rect 186998 198386 187004 198388
rect 83476 198326 187004 198386
rect 83476 198324 83482 198326
rect 186998 198324 187004 198326
rect 187068 198324 187074 198388
rect 67214 198188 67220 198252
rect 67284 198250 67290 198252
rect 67541 198250 67607 198253
rect 67284 198248 67607 198250
rect 67284 198192 67546 198248
rect 67602 198192 67607 198248
rect 67284 198190 67607 198192
rect 67284 198188 67290 198190
rect 67541 198187 67607 198190
rect 74206 198188 74212 198252
rect 74276 198250 74282 198252
rect 74349 198250 74415 198253
rect 83641 198252 83707 198253
rect 83590 198250 83596 198252
rect 74276 198248 74415 198250
rect 74276 198192 74354 198248
rect 74410 198192 74415 198248
rect 74276 198190 74415 198192
rect 83550 198190 83596 198250
rect 83660 198248 83707 198252
rect 83702 198192 83707 198248
rect 74276 198188 74282 198190
rect 74349 198187 74415 198190
rect 83590 198188 83596 198190
rect 83660 198188 83707 198192
rect 93894 198188 93900 198252
rect 93964 198250 93970 198252
rect 187550 198250 187556 198252
rect 93964 198190 187556 198250
rect 93964 198188 93970 198190
rect 187550 198188 187556 198190
rect 187620 198188 187626 198252
rect 83641 198187 83707 198188
rect 95366 198052 95372 198116
rect 95436 198114 95442 198116
rect 186814 198114 186820 198116
rect 95436 198054 186820 198114
rect 95436 198052 95442 198054
rect 186814 198052 186820 198054
rect 186884 198052 186890 198116
rect 69657 197980 69723 197981
rect 107009 197980 107075 197981
rect 69606 197978 69612 197980
rect 69566 197918 69612 197978
rect 69676 197976 69723 197980
rect 106958 197978 106964 197980
rect 69718 197920 69723 197976
rect 69606 197916 69612 197918
rect 69676 197916 69723 197920
rect 106918 197918 106964 197978
rect 107028 197976 107075 197980
rect 107070 197920 107075 197976
rect 106958 197916 106964 197918
rect 107028 197916 107075 197920
rect 108062 197916 108068 197980
rect 108132 197978 108138 197980
rect 108573 197978 108639 197981
rect 109217 197980 109283 197981
rect 109166 197978 109172 197980
rect 108132 197976 108639 197978
rect 108132 197920 108578 197976
rect 108634 197920 108639 197976
rect 108132 197918 108639 197920
rect 109126 197918 109172 197978
rect 109236 197976 109283 197980
rect 109278 197920 109283 197976
rect 108132 197916 108138 197918
rect 69657 197915 69723 197916
rect 107009 197915 107075 197916
rect 108573 197915 108639 197918
rect 109166 197916 109172 197918
rect 109236 197916 109283 197920
rect 130878 197916 130884 197980
rect 130948 197978 130954 197980
rect 188470 197978 188476 197980
rect 130948 197918 188476 197978
rect 130948 197916 130954 197918
rect 188470 197916 188476 197918
rect 188540 197916 188546 197980
rect 109217 197915 109283 197916
rect 138657 197844 138723 197845
rect 138606 197842 138612 197844
rect 138566 197782 138612 197842
rect 138676 197840 138723 197844
rect 138718 197784 138723 197840
rect 138606 197780 138612 197782
rect 138676 197780 138723 197784
rect 140998 197780 141004 197844
rect 141068 197842 141074 197844
rect 141233 197842 141299 197845
rect 143441 197844 143507 197845
rect 173249 197844 173315 197845
rect 143390 197842 143396 197844
rect 141068 197840 141299 197842
rect 141068 197784 141238 197840
rect 141294 197784 141299 197840
rect 141068 197782 141299 197784
rect 143350 197782 143396 197842
rect 143460 197840 143507 197844
rect 173198 197842 173204 197844
rect 143502 197784 143507 197840
rect 141068 197780 141074 197782
rect 138657 197779 138723 197780
rect 141233 197779 141299 197782
rect 143390 197780 143396 197782
rect 143460 197780 143507 197784
rect 173158 197782 173204 197842
rect 173268 197840 173315 197844
rect 173310 197784 173315 197840
rect 173198 197780 173204 197782
rect 173268 197780 173315 197784
rect 143441 197779 143507 197780
rect 173249 197779 173315 197780
rect 133505 197708 133571 197709
rect 148593 197708 148659 197709
rect 150985 197708 151051 197709
rect 133454 197706 133460 197708
rect 133414 197646 133460 197706
rect 133524 197704 133571 197708
rect 148542 197706 148548 197708
rect 133566 197648 133571 197704
rect 133454 197644 133460 197646
rect 133524 197644 133571 197648
rect 148502 197646 148548 197706
rect 148612 197704 148659 197708
rect 150934 197706 150940 197708
rect 148654 197648 148659 197704
rect 148542 197644 148548 197646
rect 148612 197644 148659 197648
rect 150894 197646 150940 197706
rect 151004 197704 151051 197708
rect 151046 197648 151051 197704
rect 150934 197644 150940 197646
rect 151004 197644 151051 197648
rect 133505 197643 133571 197644
rect 148593 197643 148659 197644
rect 150985 197643 151051 197644
rect 237373 197706 237439 197709
rect 237373 197704 239874 197706
rect 237373 197648 237378 197704
rect 237434 197648 239874 197704
rect 237373 197646 239874 197648
rect 237373 197643 237439 197646
rect 239814 197638 239874 197646
rect 239814 197578 240212 197638
rect 91502 197508 91508 197572
rect 91572 197570 91578 197572
rect 238518 197570 238524 197572
rect 91572 197510 238524 197570
rect 91572 197508 91578 197510
rect 238518 197508 238524 197510
rect 238588 197508 238594 197572
rect 66161 197436 66227 197437
rect 66110 197434 66116 197436
rect 66070 197374 66116 197434
rect 66180 197432 66227 197436
rect 66222 197376 66227 197432
rect 66110 197372 66116 197374
rect 66180 197372 66227 197376
rect 68318 197372 68324 197436
rect 68388 197434 68394 197436
rect 68921 197434 68987 197437
rect 68388 197432 68987 197434
rect 68388 197376 68926 197432
rect 68982 197376 68987 197432
rect 68388 197374 68987 197376
rect 68388 197372 68394 197374
rect 66161 197371 66227 197372
rect 68921 197371 68987 197374
rect 78254 197372 78260 197436
rect 78324 197434 78330 197436
rect 78581 197434 78647 197437
rect 78324 197432 78647 197434
rect 78324 197376 78586 197432
rect 78642 197376 78647 197432
rect 78324 197374 78647 197376
rect 78324 197372 78330 197374
rect 78581 197371 78647 197374
rect 80830 197372 80836 197436
rect 80900 197434 80906 197436
rect 81249 197434 81315 197437
rect 155953 197436 156019 197437
rect 155902 197434 155908 197436
rect 80900 197432 81315 197434
rect 80900 197376 81254 197432
rect 81310 197376 81315 197432
rect 80900 197374 81315 197376
rect 155862 197374 155908 197434
rect 155972 197432 156019 197436
rect 156014 197376 156019 197432
rect 80900 197372 80906 197374
rect 81249 197371 81315 197374
rect 155902 197372 155908 197374
rect 155972 197372 156019 197376
rect 155953 197371 156019 197372
rect 47853 197298 47919 197301
rect 189073 197298 189139 197301
rect 47853 197296 189139 197298
rect 47853 197240 47858 197296
rect 47914 197240 189078 197296
rect 189134 197240 189139 197296
rect 47853 197238 189139 197240
rect 47853 197235 47919 197238
rect 189073 197235 189139 197238
rect 101254 197100 101260 197164
rect 101324 197162 101330 197164
rect 234981 197162 235047 197165
rect 101324 197160 235047 197162
rect 101324 197104 234986 197160
rect 235042 197104 235047 197160
rect 101324 197102 235047 197104
rect 101324 197100 101330 197102
rect 234981 197099 235047 197102
rect 103329 197026 103395 197029
rect 235901 197026 235967 197029
rect 103329 197024 235967 197026
rect 103329 196968 103334 197024
rect 103390 196968 235906 197024
rect 235962 196968 235967 197024
rect 103329 196966 235967 196968
rect 103329 196963 103395 196966
rect 235901 196963 235967 196966
rect 100017 196890 100083 196893
rect 232773 196890 232839 196893
rect 100017 196888 232839 196890
rect 100017 196832 100022 196888
rect 100078 196832 232778 196888
rect 232834 196832 232839 196888
rect 100017 196830 232839 196832
rect 100017 196827 100083 196830
rect 232773 196827 232839 196830
rect 102225 196754 102291 196757
rect 235165 196754 235231 196757
rect 102225 196752 235231 196754
rect 102225 196696 102230 196752
rect 102286 196696 235170 196752
rect 235226 196696 235231 196752
rect 102225 196694 235231 196696
rect 102225 196691 102291 196694
rect 235165 196691 235231 196694
rect 237373 196754 237439 196757
rect 237373 196752 239874 196754
rect 237373 196696 237378 196752
rect 237434 196696 239874 196752
rect 237373 196694 239874 196696
rect 237373 196691 237439 196694
rect 239814 196686 239874 196694
rect 239814 196626 240212 196686
rect 104433 196618 104499 196621
rect 235717 196618 235783 196621
rect 104433 196616 235783 196618
rect 104433 196560 104438 196616
rect 104494 196560 235722 196616
rect 235778 196560 235783 196616
rect 104433 196558 235783 196560
rect 104433 196555 104499 196558
rect 235717 196555 235783 196558
rect 237373 195666 237439 195669
rect 237373 195664 239874 195666
rect 237373 195608 237378 195664
rect 237434 195608 239874 195664
rect 237373 195606 239874 195608
rect 237373 195603 237439 195606
rect 239814 195598 239874 195606
rect 239814 195538 240212 195598
rect 237465 194714 237531 194717
rect 237465 194712 239874 194714
rect 237465 194656 237470 194712
rect 237526 194656 239874 194712
rect 237465 194654 239874 194656
rect 237465 194651 237531 194654
rect 239814 194646 239874 194654
rect 239814 194586 240212 194646
rect 237373 193626 237439 193629
rect 237373 193624 239874 193626
rect 237373 193568 237378 193624
rect 237434 193568 239874 193624
rect 237373 193566 239874 193568
rect 237373 193563 237439 193566
rect 239814 193558 239874 193566
rect 239814 193498 240212 193558
rect 237373 192674 237439 192677
rect 237373 192672 239874 192674
rect 237373 192616 237378 192672
rect 237434 192616 239874 192672
rect 237373 192614 239874 192616
rect 237373 192611 237439 192614
rect 239814 192606 239874 192614
rect 239814 192546 240212 192606
rect 580073 192538 580139 192541
rect 583520 192538 584960 192628
rect 580073 192536 584960 192538
rect 580073 192480 580078 192536
rect 580134 192480 584960 192536
rect 580073 192478 584960 192480
rect 580073 192475 580139 192478
rect 583520 192388 584960 192478
rect 237373 191586 237439 191589
rect 237373 191584 239874 191586
rect 237373 191528 237378 191584
rect 237434 191528 239874 191584
rect 237373 191526 239874 191528
rect 237373 191523 237439 191526
rect 239814 191518 239874 191526
rect 239814 191458 240212 191518
rect 237465 190634 237531 190637
rect 237465 190632 239874 190634
rect 237465 190576 237470 190632
rect 237526 190576 239874 190632
rect 237465 190574 239874 190576
rect 237465 190571 237531 190574
rect 239814 190566 239874 190574
rect 239814 190506 240212 190566
rect 237373 189682 237439 189685
rect 237373 189680 239874 189682
rect 237373 189624 237378 189680
rect 237434 189624 239874 189680
rect 237373 189622 239874 189624
rect 237373 189619 237439 189622
rect 239814 189614 239874 189622
rect 239814 189554 240212 189614
rect -960 188866 480 188956
rect 3325 188866 3391 188869
rect -960 188864 3391 188866
rect -960 188808 3330 188864
rect 3386 188808 3391 188864
rect -960 188806 3391 188808
rect -960 188716 480 188806
rect 3325 188803 3391 188806
rect 238385 188594 238451 188597
rect 238385 188592 239874 188594
rect 238385 188536 238390 188592
rect 238446 188536 239874 188592
rect 238385 188534 239874 188536
rect 238385 188531 238451 188534
rect 239814 188526 239874 188534
rect 239814 188466 240212 188526
rect 238385 187642 238451 187645
rect 238385 187640 239874 187642
rect 238385 187584 238390 187640
rect 238446 187584 239874 187640
rect 238385 187582 239874 187584
rect 238385 187579 238451 187582
rect 239814 187574 239874 187582
rect 239814 187514 240212 187574
rect 238753 186554 238819 186557
rect 238753 186552 239874 186554
rect 238753 186496 238758 186552
rect 238814 186496 239874 186552
rect 238753 186494 239874 186496
rect 238753 186491 238819 186494
rect 239814 186486 239874 186494
rect 239814 186426 240212 186486
rect 238017 185602 238083 185605
rect 238017 185600 239874 185602
rect 238017 185544 238022 185600
rect 238078 185544 239874 185600
rect 238017 185542 239874 185544
rect 238017 185539 238083 185542
rect 239814 185534 239874 185542
rect 239814 185474 240212 185534
rect 238753 184514 238819 184517
rect 238753 184512 239874 184514
rect 238753 184456 238758 184512
rect 238814 184456 239874 184512
rect 238753 184454 239874 184456
rect 238753 184451 238819 184454
rect 239814 184446 239874 184454
rect 239814 184386 240212 184446
rect 239814 183468 240242 183528
rect 238385 183426 238451 183429
rect 239814 183426 239874 183468
rect 240182 183464 240242 183468
rect 238385 183424 239874 183426
rect 238385 183368 238390 183424
rect 238446 183368 239874 183424
rect 238385 183366 239874 183368
rect 238385 183363 238451 183366
rect 238293 182474 238359 182477
rect 238293 182472 239874 182474
rect 238293 182416 238298 182472
rect 238354 182416 239874 182472
rect 238293 182414 239874 182416
rect 238293 182411 238359 182414
rect 239814 182406 239874 182414
rect 239814 182346 240212 182406
rect 239397 181522 239463 181525
rect 239397 181520 239874 181522
rect 239397 181464 239402 181520
rect 239458 181488 239874 181520
rect 239458 181464 240242 181488
rect 239397 181462 240242 181464
rect 239397 181459 239463 181462
rect 239814 181428 240242 181462
rect 240182 181424 240242 181428
rect 238569 180570 238635 180573
rect 238569 180568 239874 180570
rect 238569 180512 238574 180568
rect 238630 180512 239874 180568
rect 238569 180510 239874 180512
rect 238569 180507 238635 180510
rect 239814 180502 239874 180510
rect 239814 180442 240212 180502
rect 370313 179754 370379 179757
rect 536782 179754 536788 179756
rect 370313 179752 536788 179754
rect 370313 179696 370318 179752
rect 370374 179696 536788 179752
rect 370313 179694 536788 179696
rect 370313 179691 370379 179694
rect 536782 179692 536788 179694
rect 536852 179692 536858 179756
rect 237966 179556 237972 179620
rect 238036 179618 238042 179620
rect 429561 179618 429627 179621
rect 238036 179616 429627 179618
rect 238036 179560 429566 179616
rect 429622 179560 429627 179616
rect 238036 179558 429627 179560
rect 238036 179556 238042 179558
rect 429561 179555 429627 179558
rect 346209 179482 346275 179485
rect 580574 179482 580580 179484
rect 346209 179480 580580 179482
rect 346209 179424 346214 179480
rect 346270 179424 580580 179480
rect 346209 179422 580580 179424
rect 346209 179419 346275 179422
rect 580574 179420 580580 179422
rect 580644 179420 580650 179484
rect 239765 179346 239831 179349
rect 469581 179346 469647 179349
rect 239765 179344 469647 179346
rect 239765 179288 239770 179344
rect 239826 179288 469586 179344
rect 469642 179288 469647 179344
rect 239765 179286 469647 179288
rect 239765 179283 239831 179286
rect 469581 179283 469647 179286
rect 239581 179210 239647 179213
rect 453573 179210 453639 179213
rect 239581 179208 453639 179210
rect 239581 179152 239586 179208
rect 239642 179152 453578 179208
rect 453634 179152 453639 179208
rect 239581 179150 453639 179152
rect 239581 179147 239647 179150
rect 453573 179147 453639 179150
rect 580165 179210 580231 179213
rect 583520 179210 584960 179300
rect 580165 179208 584960 179210
rect 580165 179152 580170 179208
rect 580226 179152 584960 179208
rect 580165 179150 584960 179152
rect 580165 179147 580231 179150
rect 373717 179074 373783 179077
rect 580206 179074 580212 179076
rect 373717 179072 580212 179074
rect 373717 179016 373722 179072
rect 373778 179016 580212 179072
rect 373717 179014 580212 179016
rect 373717 179011 373783 179014
rect 580206 179012 580212 179014
rect 580276 179012 580282 179076
rect 583520 179060 584960 179150
rect 239254 178876 239260 178940
rect 239324 178938 239330 178940
rect 445753 178938 445819 178941
rect 239324 178936 445819 178938
rect 239324 178880 445758 178936
rect 445814 178880 445819 178936
rect 239324 178878 445819 178880
rect 239324 178876 239330 178878
rect 445753 178875 445819 178878
rect 239305 178802 239371 178805
rect 437565 178802 437631 178805
rect 239305 178800 437631 178802
rect 239305 178744 239310 178800
rect 239366 178744 437570 178800
rect 437626 178744 437631 178800
rect 239305 178742 437631 178744
rect 239305 178739 239371 178742
rect 437565 178739 437631 178742
rect 449893 178666 449959 178669
rect 580390 178666 580396 178668
rect 449893 178664 580396 178666
rect 449893 178608 449898 178664
rect 449954 178608 580396 178664
rect 449893 178606 580396 178608
rect 449893 178603 449959 178606
rect 580390 178604 580396 178606
rect 580460 178604 580466 178668
rect 3601 177986 3667 177989
rect 465533 177986 465599 177989
rect 3601 177984 465599 177986
rect 3601 177928 3606 177984
rect 3662 177928 465538 177984
rect 465594 177928 465599 177984
rect 3601 177926 465599 177928
rect 3601 177923 3667 177926
rect 465533 177923 465599 177926
rect 3417 177850 3483 177853
rect 433609 177850 433675 177853
rect 3417 177848 433675 177850
rect 3417 177792 3422 177848
rect 3478 177792 433614 177848
rect 433670 177792 433675 177848
rect 3417 177790 433675 177792
rect 3417 177787 3483 177790
rect 433609 177787 433675 177790
rect 201493 177714 201559 177717
rect 421557 177714 421623 177717
rect 201493 177712 421623 177714
rect 201493 177656 201498 177712
rect 201554 177656 421562 177712
rect 421618 177656 421623 177712
rect 201493 177654 421623 177656
rect 201493 177651 201559 177654
rect 421557 177651 421623 177654
rect 218053 177578 218119 177581
rect 401409 177578 401475 177581
rect 218053 177576 401475 177578
rect 218053 177520 218058 177576
rect 218114 177520 401414 177576
rect 401470 177520 401475 177576
rect 218053 177518 401475 177520
rect 218053 177515 218119 177518
rect 401409 177515 401475 177518
rect 401593 177578 401659 177581
rect 473537 177578 473603 177581
rect 401593 177576 473603 177578
rect 401593 177520 401598 177576
rect 401654 177520 473542 177576
rect 473598 177520 473603 177576
rect 401593 177518 473603 177520
rect 401593 177515 401659 177518
rect 473537 177515 473603 177518
rect 354305 177442 354371 177445
rect 449893 177442 449959 177445
rect 354305 177440 449959 177442
rect 354305 177384 354310 177440
rect 354366 177384 449898 177440
rect 449954 177384 449959 177440
rect 354305 177382 449959 177384
rect 354305 177379 354371 177382
rect 449893 177379 449959 177382
rect 235390 176564 235396 176628
rect 235460 176626 235466 176628
rect 441705 176626 441771 176629
rect 235460 176624 441771 176626
rect 235460 176568 441710 176624
rect 441766 176568 441771 176624
rect 235460 176566 441771 176568
rect 235460 176564 235466 176566
rect 441705 176563 441771 176566
rect 235206 176428 235212 176492
rect 235276 176490 235282 176492
rect 417601 176490 417667 176493
rect 235276 176488 417667 176490
rect 235276 176432 417606 176488
rect 417662 176432 417667 176488
rect 235276 176430 417667 176432
rect 235276 176428 235282 176430
rect 417601 176427 417667 176430
rect -960 175796 480 176036
rect 583520 165732 584960 165972
rect -960 162740 480 162980
rect 580165 152690 580231 152693
rect 583520 152690 584960 152780
rect 580165 152688 584960 152690
rect 580165 152632 580170 152688
rect 580226 152632 584960 152688
rect 580165 152630 584960 152632
rect 580165 152627 580231 152630
rect 583520 152540 584960 152630
rect -960 149834 480 149924
rect 3417 149834 3483 149837
rect -960 149832 3483 149834
rect -960 149776 3422 149832
rect 3478 149776 3483 149832
rect -960 149774 3483 149776
rect -960 149684 480 149774
rect 3417 149771 3483 149774
rect 580165 139362 580231 139365
rect 583520 139362 584960 139452
rect 580165 139360 584960 139362
rect 580165 139304 580170 139360
rect 580226 139304 584960 139360
rect 580165 139302 584960 139304
rect 580165 139299 580231 139302
rect 583520 139212 584960 139302
rect -960 136778 480 136868
rect 3233 136778 3299 136781
rect -960 136776 3299 136778
rect -960 136720 3238 136776
rect 3294 136720 3299 136776
rect -960 136718 3299 136720
rect -960 136628 480 136718
rect 3233 136715 3299 136718
rect 583520 125884 584960 126124
rect -960 123572 480 123812
rect 579797 112842 579863 112845
rect 583520 112842 584960 112932
rect 579797 112840 584960 112842
rect 579797 112784 579802 112840
rect 579858 112784 584960 112840
rect 579797 112782 584960 112784
rect 579797 112779 579863 112782
rect 583520 112692 584960 112782
rect -960 110516 480 110756
rect 580165 99514 580231 99517
rect 583520 99514 584960 99604
rect 580165 99512 584960 99514
rect 580165 99456 580170 99512
rect 580226 99456 584960 99512
rect 580165 99454 584960 99456
rect 580165 99451 580231 99454
rect 583520 99364 584960 99454
rect -960 97460 480 97700
rect 583520 86036 584960 86276
rect -960 84690 480 84780
rect 3141 84690 3207 84693
rect -960 84688 3207 84690
rect -960 84632 3146 84688
rect 3202 84632 3207 84688
rect -960 84630 3207 84632
rect -960 84540 480 84630
rect 3141 84627 3207 84630
rect 580165 72994 580231 72997
rect 583520 72994 584960 73084
rect 580165 72992 584960 72994
rect 580165 72936 580170 72992
rect 580226 72936 584960 72992
rect 580165 72934 584960 72936
rect 580165 72931 580231 72934
rect 583520 72844 584960 72934
rect -960 71484 480 71724
rect 580165 59666 580231 59669
rect 583520 59666 584960 59756
rect 580165 59664 584960 59666
rect 580165 59608 580170 59664
rect 580226 59608 584960 59664
rect 580165 59606 584960 59608
rect 580165 59603 580231 59606
rect 583520 59516 584960 59606
rect -960 58428 480 58668
rect 583520 46188 584960 46428
rect -960 45522 480 45612
rect 3417 45522 3483 45525
rect -960 45520 3483 45522
rect -960 45464 3422 45520
rect 3478 45464 3483 45520
rect -960 45462 3483 45464
rect -960 45372 480 45462
rect 3417 45459 3483 45462
rect 580165 33146 580231 33149
rect 583520 33146 584960 33236
rect 580165 33144 584960 33146
rect 580165 33088 580170 33144
rect 580226 33088 584960 33144
rect 580165 33086 584960 33088
rect 580165 33083 580231 33086
rect 583520 32996 584960 33086
rect -960 32316 480 32556
rect 583520 19668 584960 19908
rect -960 19260 480 19500
rect 580165 6626 580231 6629
rect 583520 6626 584960 6716
rect 580165 6624 584960 6626
rect -960 6490 480 6580
rect 580165 6568 580170 6624
rect 580226 6568 584960 6624
rect 580165 6566 584960 6568
rect 580165 6563 580231 6566
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect 583520 6476 584960 6566
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
<< via3 >>
rect 237972 700572 238036 700636
rect 235212 700436 235276 700500
rect 239260 700300 239324 700364
rect 580212 697172 580276 697236
rect 580396 683844 580460 683908
rect 580580 630804 580644 630868
rect 235396 618292 235460 618356
rect 536788 596804 536852 596868
rect 156092 466380 156156 466444
rect 151124 466244 151188 466308
rect 81020 465564 81084 465628
rect 86172 465428 86236 465492
rect 78812 465292 78876 465356
rect 188292 465292 188356 465356
rect 91140 465216 91204 465220
rect 91140 465160 91190 465216
rect 91190 465160 91204 465216
rect 91140 465156 91204 465160
rect 93532 465156 93596 465220
rect 96108 465216 96172 465220
rect 96108 465160 96158 465216
rect 96158 465160 96172 465216
rect 96108 465156 96172 465160
rect 101260 465216 101324 465220
rect 101260 465160 101310 465216
rect 101310 465160 101324 465216
rect 101260 465156 101324 465160
rect 103652 465216 103716 465220
rect 103652 465160 103702 465216
rect 103702 465160 103716 465216
rect 103652 465156 103716 465160
rect 106228 465216 106292 465220
rect 106228 465160 106242 465216
rect 106242 465160 106292 465216
rect 106228 465156 106292 465160
rect 108436 465216 108500 465220
rect 108436 465160 108486 465216
rect 108486 465160 108500 465216
rect 108436 465156 108500 465160
rect 111012 465216 111076 465220
rect 111012 465160 111062 465216
rect 111062 465160 111076 465216
rect 111012 465156 111076 465160
rect 128676 465216 128740 465220
rect 128676 465160 128726 465216
rect 128726 465160 128740 465216
rect 128676 465156 128740 465160
rect 136036 465216 136100 465220
rect 136036 465160 136086 465216
rect 136086 465160 136100 465216
rect 136036 465156 136100 465160
rect 141004 465216 141068 465220
rect 141004 465160 141054 465216
rect 141054 465160 141068 465216
rect 141004 465156 141068 465160
rect 145972 465216 146036 465220
rect 145972 465160 146022 465216
rect 146022 465160 146036 465216
rect 145972 465156 146036 465160
rect 153332 465156 153396 465220
rect 168420 465216 168484 465220
rect 168420 465160 168470 465216
rect 168470 465160 168484 465216
rect 168420 465156 168484 465160
rect 169708 465216 169772 465220
rect 169708 465160 169758 465216
rect 169758 465160 169772 465216
rect 169708 465156 169772 465160
rect 180932 465156 180996 465220
rect 187740 465156 187804 465220
rect 131068 463992 131132 463996
rect 131068 463936 131118 463992
rect 131118 463936 131132 463992
rect 131068 463932 131132 463936
rect 83462 463720 83526 463724
rect 83462 463664 83518 463720
rect 83518 463664 83526 463720
rect 83462 463660 83526 463664
rect 88494 463720 88558 463724
rect 88494 463664 88522 463720
rect 88522 463664 88558 463720
rect 88494 463660 88558 463664
rect 98558 463720 98622 463724
rect 98558 463664 98606 463720
rect 98606 463664 98622 463720
rect 98558 463660 98622 463664
rect 113654 463720 113718 463724
rect 113654 463664 113694 463720
rect 113694 463664 113718 463720
rect 113654 463660 113718 463664
rect 116102 463720 116166 463724
rect 116102 463664 116122 463720
rect 116122 463664 116166 463720
rect 116102 463660 116166 463664
rect 118550 463720 118614 463724
rect 118550 463664 118606 463720
rect 118606 463664 118614 463720
rect 118550 463660 118614 463664
rect 120998 463720 121062 463724
rect 120998 463664 121054 463720
rect 121054 463664 121062 463720
rect 120998 463660 121062 463664
rect 123582 463720 123646 463724
rect 123582 463664 123630 463720
rect 123630 463664 123646 463720
rect 123582 463660 123646 463664
rect 125894 463660 125958 463724
rect 133510 463720 133574 463724
rect 133510 463664 133566 463720
rect 133566 463664 133574 463720
rect 133510 463660 133574 463664
rect 138406 463660 138470 463724
rect 143574 463720 143638 463724
rect 143574 463664 143630 463720
rect 143630 463664 143638 463720
rect 143574 463660 143638 463664
rect 148470 463720 148534 463724
rect 148470 463664 148506 463720
rect 148506 463664 148534 463720
rect 148470 463660 148534 463664
rect 186820 460940 186884 461004
rect 238156 456860 238220 456924
rect 238340 451420 238404 451484
rect 110934 379672 110998 379676
rect 110934 379616 110970 379672
rect 110970 379616 110998 379672
rect 110934 379612 110998 379616
rect 113518 379672 113582 379676
rect 113518 379616 113546 379672
rect 113546 379616 113582 379672
rect 113518 379612 113582 379616
rect 118278 379672 118342 379676
rect 118278 379616 118330 379672
rect 118330 379616 118342 379672
rect 118278 379612 118342 379616
rect 120998 379672 121062 379676
rect 120998 379616 121054 379672
rect 121054 379616 121062 379672
rect 120998 379612 121062 379616
rect 123446 379672 123510 379676
rect 123446 379616 123482 379672
rect 123482 379616 123510 379672
rect 123446 379612 123510 379616
rect 130926 379672 130990 379676
rect 130926 379616 130934 379672
rect 130934 379616 130990 379672
rect 130926 379612 130990 379616
rect 143438 379612 143502 379676
rect 86998 379536 87062 379540
rect 86998 379480 87050 379536
rect 87050 379480 87062 379536
rect 86998 379476 87062 379480
rect 88086 379476 88150 379540
rect 89446 379536 89510 379540
rect 89446 379480 89498 379536
rect 89498 379480 89510 379536
rect 89446 379476 89510 379480
rect 90670 379536 90734 379540
rect 90670 379480 90730 379536
rect 90730 379480 90734 379536
rect 90670 379476 90734 379480
rect 115980 379536 116044 379540
rect 115980 379480 116030 379536
rect 116030 379480 116044 379536
rect 115980 379476 116044 379480
rect 150940 379536 151004 379540
rect 150940 379480 150990 379536
rect 150990 379480 151004 379536
rect 150940 379476 151004 379480
rect 101260 379340 101324 379404
rect 103284 379204 103348 379268
rect 238340 379204 238404 379268
rect 109172 379068 109236 379132
rect 98684 378932 98748 378996
rect 67220 378116 67284 378180
rect 74212 378116 74276 378180
rect 77708 378116 77772 378180
rect 81204 378116 81268 378180
rect 91876 378116 91940 378180
rect 95924 378116 95988 378180
rect 99788 378116 99852 378180
rect 103652 378116 103716 378180
rect 128492 378116 128556 378180
rect 145972 378116 146036 378180
rect 153332 378116 153396 378180
rect 85804 377980 85868 378044
rect 92796 378040 92860 378044
rect 92796 377984 92846 378040
rect 92846 377984 92860 378040
rect 92796 377980 92860 377984
rect 93900 378040 93964 378044
rect 93900 377984 93950 378040
rect 93950 377984 93964 378040
rect 93900 377980 93964 377984
rect 95188 378040 95252 378044
rect 95188 377984 95238 378040
rect 95238 377984 95252 378040
rect 95188 377980 95252 377984
rect 97580 378040 97644 378044
rect 97580 377984 97630 378040
rect 97630 377984 97644 378040
rect 97580 377980 97644 377984
rect 106044 378040 106108 378044
rect 106044 377984 106094 378040
rect 106094 377984 106108 378040
rect 106044 377980 106108 377984
rect 108436 378040 108500 378044
rect 108436 377984 108486 378040
rect 108486 377984 108500 378040
rect 108436 377980 108500 377984
rect 125916 378040 125980 378044
rect 125916 377984 125966 378040
rect 125966 377984 125980 378040
rect 125916 377980 125980 377984
rect 133460 378040 133524 378044
rect 133460 377984 133510 378040
rect 133510 377984 133524 378040
rect 133460 377980 133524 377984
rect 136036 378040 136100 378044
rect 136036 377984 136086 378040
rect 136086 377984 136100 378040
rect 136036 377980 136100 377984
rect 138612 378040 138676 378044
rect 138612 377984 138662 378040
rect 138662 377984 138676 378040
rect 138612 377980 138676 377984
rect 141004 377980 141068 378044
rect 148548 378040 148612 378044
rect 148548 377984 148598 378040
rect 148598 377984 148612 378040
rect 148548 377980 148612 377984
rect 155908 378040 155972 378044
rect 155908 377984 155958 378040
rect 155958 377984 155972 378040
rect 155908 377980 155972 377984
rect 96476 377904 96540 377908
rect 96476 377848 96490 377904
rect 96490 377848 96540 377904
rect 96476 377844 96540 377848
rect 104388 377844 104452 377908
rect 238156 377844 238220 377908
rect 101076 377708 101140 377772
rect 106964 377708 107028 377772
rect 108068 377572 108132 377636
rect 105860 377436 105924 377500
rect 186820 377436 186884 377500
rect 187740 377300 187804 377364
rect 173204 377164 173268 377228
rect 66116 377088 66180 377092
rect 66116 377032 66166 377088
rect 66166 377032 66180 377088
rect 66116 377028 66180 377032
rect 68324 377028 68388 377092
rect 69612 377028 69676 377092
rect 70532 377028 70596 377092
rect 71820 377028 71884 377092
rect 75500 377028 75564 377092
rect 76604 377028 76668 377092
rect 78260 377088 78324 377092
rect 78260 377032 78310 377088
rect 78310 377032 78324 377088
rect 78260 377028 78324 377032
rect 78812 377028 78876 377092
rect 80100 377028 80164 377092
rect 82492 377028 82556 377092
rect 83596 377028 83660 377092
rect 84516 377028 84580 377092
rect 85988 377028 86052 377092
rect 88564 377028 88628 377092
rect 91140 377028 91204 377092
rect 93532 377028 93596 377092
rect 98316 377028 98380 377092
rect 102180 377028 102244 377092
rect 73108 376892 73172 376956
rect 80836 376892 80900 376956
rect 83412 376892 83476 376956
rect 173388 376892 173452 376956
rect 188292 317460 188356 317524
rect 116164 286452 116228 286516
rect 136036 286316 136100 286380
rect 169708 286316 169772 286380
rect 168420 286180 168484 286244
rect 125916 286044 125980 286108
rect 131068 286044 131132 286108
rect 133460 286044 133524 286108
rect 108436 285908 108500 285972
rect 111012 285908 111076 285972
rect 78812 285636 78876 285700
rect 81020 285636 81084 285700
rect 83412 285636 83476 285700
rect 188292 285772 188356 285836
rect 86172 285636 86236 285700
rect 88564 285636 88628 285700
rect 93532 285636 93596 285700
rect 101260 285636 101324 285700
rect 103836 285636 103900 285700
rect 106228 285696 106292 285700
rect 106228 285640 106242 285696
rect 106242 285640 106292 285696
rect 106228 285636 106292 285640
rect 120764 285636 120828 285700
rect 138428 285636 138492 285700
rect 141004 285636 141068 285700
rect 143580 285636 143644 285700
rect 145604 285636 145668 285700
rect 148548 285636 148612 285700
rect 151124 285636 151188 285700
rect 154068 285636 154132 285700
rect 156092 285636 156156 285700
rect 96108 285152 96172 285156
rect 96108 285096 96158 285152
rect 96158 285096 96172 285152
rect 96108 285092 96172 285096
rect 113772 285152 113836 285156
rect 113772 285096 113822 285152
rect 113822 285096 113836 285152
rect 113772 285092 113836 285096
rect 123524 285152 123588 285156
rect 123524 285096 123574 285152
rect 123574 285096 123588 285152
rect 123524 285092 123588 285096
rect 128676 285152 128740 285156
rect 128676 285096 128726 285152
rect 128726 285096 128740 285152
rect 128676 285092 128740 285096
rect 98500 285016 98564 285020
rect 98500 284960 98550 285016
rect 98550 284960 98564 285016
rect 98500 284956 98564 284960
rect 118556 285016 118620 285020
rect 118556 284960 118606 285016
rect 118606 284960 118620 285016
rect 118556 284956 118620 284960
rect 91140 284880 91204 284884
rect 91140 284824 91190 284880
rect 91190 284824 91204 284880
rect 91140 284820 91204 284824
rect 180748 284064 180812 284068
rect 180748 284008 180762 284064
rect 180762 284008 180812 284064
rect 180748 284004 180812 284008
rect 238156 277612 238220 277676
rect 186820 270540 186884 270604
rect 238340 268500 238404 268564
rect 238524 262380 238588 262444
rect 187004 234636 187068 234700
rect 188476 222804 188540 222868
rect 187556 200636 187620 200700
rect 238340 200772 238404 200836
rect 70532 199472 70596 199476
rect 70532 199416 70582 199472
rect 70582 199416 70596 199472
rect 70532 199412 70596 199416
rect 77708 199472 77772 199476
rect 77708 199416 77758 199472
rect 77758 199416 77772 199472
rect 77708 199412 77772 199416
rect 78812 199472 78876 199476
rect 78812 199416 78862 199472
rect 78862 199416 78876 199472
rect 78812 199412 78876 199416
rect 88564 199472 88628 199476
rect 88564 199416 88614 199472
rect 88614 199416 88628 199472
rect 88564 199412 88628 199416
rect 91140 199472 91204 199476
rect 91140 199416 91190 199472
rect 91190 199416 91204 199472
rect 91140 199412 91204 199416
rect 103652 199472 103716 199476
rect 103652 199416 103702 199472
rect 103702 199416 103716 199472
rect 103652 199412 103716 199416
rect 111012 199472 111076 199476
rect 111012 199416 111062 199472
rect 111062 199416 111076 199472
rect 111012 199412 111076 199416
rect 188292 199140 188356 199204
rect 98684 199004 98748 199068
rect 96476 198868 96540 198932
rect 136036 198732 136100 198796
rect 71820 198656 71884 198660
rect 71820 198600 71870 198656
rect 71870 198600 71884 198656
rect 71820 198596 71884 198600
rect 75500 198656 75564 198660
rect 75500 198600 75550 198656
rect 75550 198600 75564 198656
rect 75500 198596 75564 198600
rect 76604 198596 76668 198660
rect 80100 198656 80164 198660
rect 80100 198600 80150 198656
rect 80150 198600 80164 198656
rect 80100 198596 80164 198600
rect 81388 198656 81452 198660
rect 81388 198600 81402 198656
rect 81402 198600 81452 198656
rect 81388 198596 81452 198600
rect 82492 198656 82556 198660
rect 82492 198600 82542 198656
rect 82542 198600 82556 198656
rect 82492 198596 82556 198600
rect 84516 198656 84580 198660
rect 84516 198600 84566 198656
rect 84566 198600 84580 198656
rect 84516 198596 84580 198600
rect 86172 198656 86236 198660
rect 86172 198600 86222 198656
rect 86222 198600 86236 198656
rect 86172 198596 86236 198600
rect 87092 198596 87156 198660
rect 92796 198656 92860 198660
rect 92796 198600 92846 198656
rect 92846 198600 92860 198656
rect 92796 198596 92860 198600
rect 93532 198656 93596 198660
rect 93532 198600 93582 198656
rect 93582 198600 93596 198656
rect 93532 198596 93596 198600
rect 95924 198656 95988 198660
rect 95924 198600 95974 198656
rect 95974 198600 95988 198656
rect 95924 198596 95988 198600
rect 97580 198596 97644 198660
rect 104388 198656 104452 198660
rect 104388 198600 104438 198656
rect 104438 198600 104452 198656
rect 85804 198520 85868 198524
rect 85804 198464 85854 198520
rect 85854 198464 85868 198520
rect 85804 198460 85868 198464
rect 88196 198520 88260 198524
rect 88196 198464 88246 198520
rect 88246 198464 88260 198520
rect 88196 198460 88260 198464
rect 89484 198520 89548 198524
rect 89484 198464 89534 198520
rect 89534 198464 89548 198520
rect 89484 198460 89548 198464
rect 90772 198520 90836 198524
rect 90772 198464 90822 198520
rect 90822 198464 90836 198520
rect 90772 198460 90836 198464
rect 98316 198520 98380 198524
rect 98316 198464 98366 198520
rect 98366 198464 98380 198520
rect 98316 198460 98380 198464
rect 99788 198460 99852 198524
rect 100892 198520 100956 198524
rect 100892 198464 100942 198520
rect 100942 198464 100956 198520
rect 100892 198460 100956 198464
rect 102180 198520 102244 198524
rect 102180 198464 102230 198520
rect 102230 198464 102244 198520
rect 102180 198460 102244 198464
rect 103284 198520 103348 198524
rect 103284 198464 103334 198520
rect 103334 198464 103348 198520
rect 103284 198460 103348 198464
rect 104388 198596 104452 198600
rect 105860 198656 105924 198660
rect 105860 198600 105910 198656
rect 105910 198600 105924 198656
rect 105860 198596 105924 198600
rect 106044 198656 106108 198660
rect 106044 198600 106094 198656
rect 106094 198600 106108 198656
rect 106044 198596 106108 198600
rect 108436 198656 108500 198660
rect 108436 198600 108486 198656
rect 108486 198600 108500 198656
rect 108436 198596 108500 198600
rect 113588 198656 113652 198660
rect 113588 198600 113638 198656
rect 113638 198600 113652 198656
rect 113588 198596 113652 198600
rect 115980 198596 116044 198660
rect 118372 198656 118436 198660
rect 118372 198600 118422 198656
rect 118422 198600 118436 198656
rect 118372 198596 118436 198600
rect 120948 198656 121012 198660
rect 120948 198600 120998 198656
rect 120998 198600 121012 198656
rect 120948 198596 121012 198600
rect 123524 198656 123588 198660
rect 123524 198600 123574 198656
rect 123574 198600 123588 198656
rect 123524 198596 123588 198600
rect 125916 198596 125980 198660
rect 128492 198596 128556 198660
rect 145972 198656 146036 198660
rect 145972 198600 146022 198656
rect 146022 198600 146036 198656
rect 145972 198596 146036 198600
rect 153332 198656 153396 198660
rect 153332 198600 153382 198656
rect 153382 198600 153396 198656
rect 153332 198596 153396 198600
rect 173388 198656 173452 198660
rect 173388 198600 173438 198656
rect 173438 198600 173452 198656
rect 173388 198596 173452 198600
rect 238156 198460 238220 198524
rect 73108 198324 73172 198388
rect 83412 198324 83476 198388
rect 187004 198324 187068 198388
rect 67220 198188 67284 198252
rect 74212 198188 74276 198252
rect 83596 198248 83660 198252
rect 83596 198192 83646 198248
rect 83646 198192 83660 198248
rect 83596 198188 83660 198192
rect 93900 198188 93964 198252
rect 187556 198188 187620 198252
rect 95372 198052 95436 198116
rect 186820 198052 186884 198116
rect 69612 197976 69676 197980
rect 69612 197920 69662 197976
rect 69662 197920 69676 197976
rect 69612 197916 69676 197920
rect 106964 197976 107028 197980
rect 106964 197920 107014 197976
rect 107014 197920 107028 197976
rect 106964 197916 107028 197920
rect 108068 197916 108132 197980
rect 109172 197976 109236 197980
rect 109172 197920 109222 197976
rect 109222 197920 109236 197976
rect 109172 197916 109236 197920
rect 130884 197916 130948 197980
rect 188476 197916 188540 197980
rect 138612 197840 138676 197844
rect 138612 197784 138662 197840
rect 138662 197784 138676 197840
rect 138612 197780 138676 197784
rect 141004 197780 141068 197844
rect 143396 197840 143460 197844
rect 143396 197784 143446 197840
rect 143446 197784 143460 197840
rect 143396 197780 143460 197784
rect 173204 197840 173268 197844
rect 173204 197784 173254 197840
rect 173254 197784 173268 197840
rect 173204 197780 173268 197784
rect 133460 197704 133524 197708
rect 133460 197648 133510 197704
rect 133510 197648 133524 197704
rect 133460 197644 133524 197648
rect 148548 197704 148612 197708
rect 148548 197648 148598 197704
rect 148598 197648 148612 197704
rect 148548 197644 148612 197648
rect 150940 197704 151004 197708
rect 150940 197648 150990 197704
rect 150990 197648 151004 197704
rect 150940 197644 151004 197648
rect 91508 197508 91572 197572
rect 238524 197508 238588 197572
rect 66116 197432 66180 197436
rect 66116 197376 66166 197432
rect 66166 197376 66180 197432
rect 66116 197372 66180 197376
rect 68324 197372 68388 197436
rect 78260 197372 78324 197436
rect 80836 197372 80900 197436
rect 155908 197432 155972 197436
rect 155908 197376 155958 197432
rect 155958 197376 155972 197432
rect 155908 197372 155972 197376
rect 101260 197100 101324 197164
rect 536788 179692 536852 179756
rect 237972 179556 238036 179620
rect 580580 179420 580644 179484
rect 580212 179012 580276 179076
rect 239260 178876 239324 178940
rect 580396 178604 580460 178668
rect 235396 176564 235460 176628
rect 235212 176428 235276 176492
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 680614 -8106 711002
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 -8106 680614
rect -8726 680294 -8106 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 -8106 680294
rect -8726 644614 -8106 680058
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 -8106 644614
rect -8726 644294 -8106 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 -8106 644294
rect -8726 608614 -8106 644058
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 -8106 608614
rect -8726 608294 -8106 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 -8106 608294
rect -8726 572614 -8106 608058
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 -8106 572614
rect -8726 572294 -8106 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 -8106 572294
rect -8726 536614 -8106 572058
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 -8106 536614
rect -8726 536294 -8106 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 -8106 536294
rect -8726 500614 -8106 536058
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 -8106 500614
rect -8726 500294 -8106 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 -8106 500294
rect -8726 464614 -8106 500058
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 -8106 464614
rect -8726 464294 -8106 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 -8106 464294
rect -8726 428614 -8106 464058
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 -8106 428614
rect -8726 428294 -8106 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 -8106 428294
rect -8726 392614 -8106 428058
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 -8106 392614
rect -8726 392294 -8106 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 -8106 392294
rect -8726 356614 -8106 392058
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 -8106 356614
rect -8726 356294 -8106 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 -8106 356294
rect -8726 320614 -8106 356058
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 -8106 320614
rect -8726 320294 -8106 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 -8106 320294
rect -8726 284614 -8106 320058
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 -8106 284614
rect -8726 284294 -8106 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 -8106 284294
rect -8726 248614 -8106 284058
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 -8106 248614
rect -8726 248294 -8106 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 -8106 248294
rect -8726 212614 -8106 248058
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 -8106 212614
rect -8726 212294 -8106 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 -8106 212294
rect -8726 176614 -8106 212058
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 -8106 176614
rect -8726 176294 -8106 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 -8106 176294
rect -8726 140614 -8106 176058
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 -8106 140614
rect -8726 140294 -8106 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 -8106 140294
rect -8726 104614 -8106 140058
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 -8106 104614
rect -8726 104294 -8106 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 -8106 104294
rect -8726 68614 -8106 104058
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 -8106 68614
rect -8726 68294 -8106 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 -8106 68294
rect -8726 32614 -8106 68058
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 -8106 32614
rect -8726 32294 -8106 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 -8106 32294
rect -8726 -7066 -8106 32058
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 698614 -7146 710042
rect 12954 710598 13574 711590
rect 12954 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 13574 710598
rect 12954 710278 13574 710362
rect 12954 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 13574 710278
rect -7766 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 -7146 698614
rect -7766 698294 -7146 698378
rect -7766 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 -7146 698294
rect -7766 662614 -7146 698058
rect -7766 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 -7146 662614
rect -7766 662294 -7146 662378
rect -7766 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 -7146 662294
rect -7766 626614 -7146 662058
rect -7766 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 -7146 626614
rect -7766 626294 -7146 626378
rect -7766 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 -7146 626294
rect -7766 590614 -7146 626058
rect -7766 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 -7146 590614
rect -7766 590294 -7146 590378
rect -7766 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 -7146 590294
rect -7766 554614 -7146 590058
rect -7766 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 -7146 554614
rect -7766 554294 -7146 554378
rect -7766 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 -7146 554294
rect -7766 518614 -7146 554058
rect -7766 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 -7146 518614
rect -7766 518294 -7146 518378
rect -7766 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 -7146 518294
rect -7766 482614 -7146 518058
rect -7766 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 -7146 482614
rect -7766 482294 -7146 482378
rect -7766 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 -7146 482294
rect -7766 446614 -7146 482058
rect -7766 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 -7146 446614
rect -7766 446294 -7146 446378
rect -7766 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 -7146 446294
rect -7766 410614 -7146 446058
rect -7766 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 -7146 410614
rect -7766 410294 -7146 410378
rect -7766 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 -7146 410294
rect -7766 374614 -7146 410058
rect -7766 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 -7146 374614
rect -7766 374294 -7146 374378
rect -7766 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 -7146 374294
rect -7766 338614 -7146 374058
rect -7766 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 -7146 338614
rect -7766 338294 -7146 338378
rect -7766 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 -7146 338294
rect -7766 302614 -7146 338058
rect -7766 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 -7146 302614
rect -7766 302294 -7146 302378
rect -7766 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 -7146 302294
rect -7766 266614 -7146 302058
rect -7766 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 -7146 266614
rect -7766 266294 -7146 266378
rect -7766 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 -7146 266294
rect -7766 230614 -7146 266058
rect -7766 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 -7146 230614
rect -7766 230294 -7146 230378
rect -7766 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 -7146 230294
rect -7766 194614 -7146 230058
rect -7766 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 -7146 194614
rect -7766 194294 -7146 194378
rect -7766 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 -7146 194294
rect -7766 158614 -7146 194058
rect -7766 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 -7146 158614
rect -7766 158294 -7146 158378
rect -7766 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 -7146 158294
rect -7766 122614 -7146 158058
rect -7766 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 -7146 122614
rect -7766 122294 -7146 122378
rect -7766 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 -7146 122294
rect -7766 86614 -7146 122058
rect -7766 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 -7146 86614
rect -7766 86294 -7146 86378
rect -7766 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 -7146 86294
rect -7766 50614 -7146 86058
rect -7766 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 -7146 50614
rect -7766 50294 -7146 50378
rect -7766 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 -7146 50294
rect -7766 14614 -7146 50058
rect -7766 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 -7146 14614
rect -7766 14294 -7146 14378
rect -7766 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 -7146 14294
rect -7766 -6106 -7146 14058
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 676894 -6186 709082
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 -6186 676894
rect -6806 676574 -6186 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 -6186 676574
rect -6806 640894 -6186 676338
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 -6186 640894
rect -6806 640574 -6186 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 -6186 640574
rect -6806 604894 -6186 640338
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 -6186 604894
rect -6806 604574 -6186 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 -6186 604574
rect -6806 568894 -6186 604338
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 -6186 568894
rect -6806 568574 -6186 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 -6186 568574
rect -6806 532894 -6186 568338
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 -6186 532894
rect -6806 532574 -6186 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 -6186 532574
rect -6806 496894 -6186 532338
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 -6186 496894
rect -6806 496574 -6186 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 -6186 496574
rect -6806 460894 -6186 496338
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 -6186 460894
rect -6806 460574 -6186 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 -6186 460574
rect -6806 424894 -6186 460338
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 -6186 424894
rect -6806 424574 -6186 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 -6186 424574
rect -6806 388894 -6186 424338
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 -6186 388894
rect -6806 388574 -6186 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 -6186 388574
rect -6806 352894 -6186 388338
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 -6186 352894
rect -6806 352574 -6186 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 -6186 352574
rect -6806 316894 -6186 352338
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 -6186 316894
rect -6806 316574 -6186 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 -6186 316574
rect -6806 280894 -6186 316338
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 -6186 280894
rect -6806 280574 -6186 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 -6186 280574
rect -6806 244894 -6186 280338
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 -6186 244894
rect -6806 244574 -6186 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 -6186 244574
rect -6806 208894 -6186 244338
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 -6186 208894
rect -6806 208574 -6186 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 -6186 208574
rect -6806 172894 -6186 208338
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 -6186 172894
rect -6806 172574 -6186 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 -6186 172574
rect -6806 136894 -6186 172338
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 -6186 136894
rect -6806 136574 -6186 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 -6186 136574
rect -6806 100894 -6186 136338
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 -6186 100894
rect -6806 100574 -6186 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 -6186 100574
rect -6806 64894 -6186 100338
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 -6186 64894
rect -6806 64574 -6186 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 -6186 64574
rect -6806 28894 -6186 64338
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 -6186 28894
rect -6806 28574 -6186 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 -6186 28574
rect -6806 -5146 -6186 28338
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 694894 -5226 708122
rect 9234 708678 9854 709670
rect 9234 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 9854 708678
rect 9234 708358 9854 708442
rect 9234 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 9854 708358
rect -5846 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 -5226 694894
rect -5846 694574 -5226 694658
rect -5846 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 -5226 694574
rect -5846 658894 -5226 694338
rect -5846 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 -5226 658894
rect -5846 658574 -5226 658658
rect -5846 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 -5226 658574
rect -5846 622894 -5226 658338
rect -5846 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 -5226 622894
rect -5846 622574 -5226 622658
rect -5846 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 -5226 622574
rect -5846 586894 -5226 622338
rect -5846 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 -5226 586894
rect -5846 586574 -5226 586658
rect -5846 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 -5226 586574
rect -5846 550894 -5226 586338
rect -5846 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 -5226 550894
rect -5846 550574 -5226 550658
rect -5846 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 -5226 550574
rect -5846 514894 -5226 550338
rect -5846 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 -5226 514894
rect -5846 514574 -5226 514658
rect -5846 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 -5226 514574
rect -5846 478894 -5226 514338
rect -5846 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 -5226 478894
rect -5846 478574 -5226 478658
rect -5846 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 -5226 478574
rect -5846 442894 -5226 478338
rect -5846 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 -5226 442894
rect -5846 442574 -5226 442658
rect -5846 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 -5226 442574
rect -5846 406894 -5226 442338
rect -5846 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 -5226 406894
rect -5846 406574 -5226 406658
rect -5846 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 -5226 406574
rect -5846 370894 -5226 406338
rect -5846 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 -5226 370894
rect -5846 370574 -5226 370658
rect -5846 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 -5226 370574
rect -5846 334894 -5226 370338
rect -5846 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 -5226 334894
rect -5846 334574 -5226 334658
rect -5846 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 -5226 334574
rect -5846 298894 -5226 334338
rect -5846 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 -5226 298894
rect -5846 298574 -5226 298658
rect -5846 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 -5226 298574
rect -5846 262894 -5226 298338
rect -5846 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 -5226 262894
rect -5846 262574 -5226 262658
rect -5846 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 -5226 262574
rect -5846 226894 -5226 262338
rect -5846 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 -5226 226894
rect -5846 226574 -5226 226658
rect -5846 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 -5226 226574
rect -5846 190894 -5226 226338
rect -5846 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 -5226 190894
rect -5846 190574 -5226 190658
rect -5846 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 -5226 190574
rect -5846 154894 -5226 190338
rect -5846 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 -5226 154894
rect -5846 154574 -5226 154658
rect -5846 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 -5226 154574
rect -5846 118894 -5226 154338
rect -5846 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 -5226 118894
rect -5846 118574 -5226 118658
rect -5846 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 -5226 118574
rect -5846 82894 -5226 118338
rect -5846 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 -5226 82894
rect -5846 82574 -5226 82658
rect -5846 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 -5226 82574
rect -5846 46894 -5226 82338
rect -5846 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 -5226 46894
rect -5846 46574 -5226 46658
rect -5846 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 -5226 46574
rect -5846 10894 -5226 46338
rect -5846 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 -5226 10894
rect -5846 10574 -5226 10658
rect -5846 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 -5226 10574
rect -5846 -4186 -5226 10338
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 673174 -4266 707162
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 -4266 673174
rect -4886 672854 -4266 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 -4266 672854
rect -4886 637174 -4266 672618
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 -4266 637174
rect -4886 636854 -4266 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 -4266 636854
rect -4886 601174 -4266 636618
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 -4266 601174
rect -4886 600854 -4266 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 -4266 600854
rect -4886 565174 -4266 600618
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 -4266 565174
rect -4886 564854 -4266 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 -4266 564854
rect -4886 529174 -4266 564618
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 -4266 529174
rect -4886 528854 -4266 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 -4266 528854
rect -4886 493174 -4266 528618
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 -4266 493174
rect -4886 492854 -4266 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 -4266 492854
rect -4886 457174 -4266 492618
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 -4266 457174
rect -4886 456854 -4266 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 -4266 456854
rect -4886 421174 -4266 456618
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 -4266 421174
rect -4886 420854 -4266 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 -4266 420854
rect -4886 385174 -4266 420618
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 -4266 385174
rect -4886 384854 -4266 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 -4266 384854
rect -4886 349174 -4266 384618
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 -4266 349174
rect -4886 348854 -4266 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 -4266 348854
rect -4886 313174 -4266 348618
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 -4266 313174
rect -4886 312854 -4266 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 -4266 312854
rect -4886 277174 -4266 312618
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 -4266 277174
rect -4886 276854 -4266 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 -4266 276854
rect -4886 241174 -4266 276618
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 -4266 241174
rect -4886 240854 -4266 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 -4266 240854
rect -4886 205174 -4266 240618
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 -4266 205174
rect -4886 204854 -4266 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 -4266 204854
rect -4886 169174 -4266 204618
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 -4266 169174
rect -4886 168854 -4266 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 -4266 168854
rect -4886 133174 -4266 168618
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 -4266 133174
rect -4886 132854 -4266 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 -4266 132854
rect -4886 97174 -4266 132618
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 -4266 97174
rect -4886 96854 -4266 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 -4266 96854
rect -4886 61174 -4266 96618
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 -4266 61174
rect -4886 60854 -4266 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 -4266 60854
rect -4886 25174 -4266 60618
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 -4266 25174
rect -4886 24854 -4266 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 -4266 24854
rect -4886 -3226 -4266 24618
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 691174 -3306 706202
rect 5514 706758 6134 707750
rect 5514 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 6134 706758
rect 5514 706438 6134 706522
rect 5514 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 6134 706438
rect -3926 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 -3306 691174
rect -3926 690854 -3306 690938
rect -3926 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 -3306 690854
rect -3926 655174 -3306 690618
rect -3926 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 -3306 655174
rect -3926 654854 -3306 654938
rect -3926 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 -3306 654854
rect -3926 619174 -3306 654618
rect -3926 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 -3306 619174
rect -3926 618854 -3306 618938
rect -3926 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 -3306 618854
rect -3926 583174 -3306 618618
rect -3926 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 -3306 583174
rect -3926 582854 -3306 582938
rect -3926 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 -3306 582854
rect -3926 547174 -3306 582618
rect -3926 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 -3306 547174
rect -3926 546854 -3306 546938
rect -3926 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 -3306 546854
rect -3926 511174 -3306 546618
rect -3926 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 -3306 511174
rect -3926 510854 -3306 510938
rect -3926 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 -3306 510854
rect -3926 475174 -3306 510618
rect -3926 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 -3306 475174
rect -3926 474854 -3306 474938
rect -3926 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 -3306 474854
rect -3926 439174 -3306 474618
rect -3926 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 -3306 439174
rect -3926 438854 -3306 438938
rect -3926 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 -3306 438854
rect -3926 403174 -3306 438618
rect -3926 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 -3306 403174
rect -3926 402854 -3306 402938
rect -3926 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 -3306 402854
rect -3926 367174 -3306 402618
rect -3926 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 -3306 367174
rect -3926 366854 -3306 366938
rect -3926 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 -3306 366854
rect -3926 331174 -3306 366618
rect -3926 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 -3306 331174
rect -3926 330854 -3306 330938
rect -3926 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 -3306 330854
rect -3926 295174 -3306 330618
rect -3926 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 -3306 295174
rect -3926 294854 -3306 294938
rect -3926 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 -3306 294854
rect -3926 259174 -3306 294618
rect -3926 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 -3306 259174
rect -3926 258854 -3306 258938
rect -3926 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 -3306 258854
rect -3926 223174 -3306 258618
rect -3926 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 -3306 223174
rect -3926 222854 -3306 222938
rect -3926 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 -3306 222854
rect -3926 187174 -3306 222618
rect -3926 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 -3306 187174
rect -3926 186854 -3306 186938
rect -3926 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 -3306 186854
rect -3926 151174 -3306 186618
rect -3926 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 -3306 151174
rect -3926 150854 -3306 150938
rect -3926 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 -3306 150854
rect -3926 115174 -3306 150618
rect -3926 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 -3306 115174
rect -3926 114854 -3306 114938
rect -3926 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 -3306 114854
rect -3926 79174 -3306 114618
rect -3926 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 -3306 79174
rect -3926 78854 -3306 78938
rect -3926 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 -3306 78854
rect -3926 43174 -3306 78618
rect -3926 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 -3306 43174
rect -3926 42854 -3306 42938
rect -3926 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 -3306 42854
rect -3926 7174 -3306 42618
rect -3926 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 -3306 7174
rect -3926 6854 -3306 6938
rect -3926 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 -3306 6854
rect -3926 -2266 -3306 6618
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 669454 -2346 705242
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 -2346 669454
rect -2966 669134 -2346 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 -2346 669134
rect -2966 633454 -2346 668898
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 -2346 633454
rect -2966 633134 -2346 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 -2346 633134
rect -2966 597454 -2346 632898
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 -2346 597454
rect -2966 597134 -2346 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 -2346 597134
rect -2966 561454 -2346 596898
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 -2346 561454
rect -2966 561134 -2346 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 -2346 561134
rect -2966 525454 -2346 560898
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 -2346 525454
rect -2966 525134 -2346 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 -2346 525134
rect -2966 489454 -2346 524898
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 -2346 489454
rect -2966 489134 -2346 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 -2346 489134
rect -2966 453454 -2346 488898
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 -2346 453454
rect -2966 453134 -2346 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 -2346 453134
rect -2966 417454 -2346 452898
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 -2346 417454
rect -2966 417134 -2346 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 -2346 417134
rect -2966 381454 -2346 416898
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 -2346 381454
rect -2966 381134 -2346 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 -2346 381134
rect -2966 345454 -2346 380898
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 -2346 345454
rect -2966 345134 -2346 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 -2346 345134
rect -2966 309454 -2346 344898
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 -2346 309454
rect -2966 309134 -2346 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 -2346 309134
rect -2966 273454 -2346 308898
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 -2346 273454
rect -2966 273134 -2346 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 -2346 273134
rect -2966 237454 -2346 272898
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 -2346 237454
rect -2966 237134 -2346 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 -2346 237134
rect -2966 201454 -2346 236898
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 -2346 201454
rect -2966 201134 -2346 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 -2346 201134
rect -2966 165454 -2346 200898
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 -2346 165454
rect -2966 165134 -2346 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 -2346 165134
rect -2966 129454 -2346 164898
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 -2346 129454
rect -2966 129134 -2346 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 -2346 129134
rect -2966 93454 -2346 128898
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 -2346 93454
rect -2966 93134 -2346 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 -2346 93134
rect -2966 57454 -2346 92898
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 -2346 57454
rect -2966 57134 -2346 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 -2346 57134
rect -2966 21454 -2346 56898
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 -2346 21454
rect -2966 21134 -2346 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 -2346 21134
rect -2966 -1306 -2346 20898
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 705830
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 1794 -1894 2414 -902
rect 5514 691174 6134 706202
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect 5514 -2266 6134 6618
rect 5514 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 6134 -2266
rect 5514 -2586 6134 -2502
rect 5514 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 6134 -2586
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect 5514 -3814 6134 -2822
rect 9234 694894 9854 708122
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 658894 9854 694338
rect 9234 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 9854 658894
rect 9234 658574 9854 658658
rect 9234 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 9854 658574
rect 9234 622894 9854 658338
rect 9234 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 9854 622894
rect 9234 622574 9854 622658
rect 9234 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 9854 622574
rect 9234 586894 9854 622338
rect 9234 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 9854 586894
rect 9234 586574 9854 586658
rect 9234 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 9854 586574
rect 9234 550894 9854 586338
rect 9234 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 9854 550894
rect 9234 550574 9854 550658
rect 9234 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 9854 550574
rect 9234 514894 9854 550338
rect 9234 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 9854 514894
rect 9234 514574 9854 514658
rect 9234 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 9854 514574
rect 9234 478894 9854 514338
rect 9234 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 9854 478894
rect 9234 478574 9854 478658
rect 9234 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 9854 478574
rect 9234 442894 9854 478338
rect 9234 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 9854 442894
rect 9234 442574 9854 442658
rect 9234 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 9854 442574
rect 9234 406894 9854 442338
rect 9234 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 9854 406894
rect 9234 406574 9854 406658
rect 9234 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 9854 406574
rect 9234 370894 9854 406338
rect 9234 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 9854 370894
rect 9234 370574 9854 370658
rect 9234 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 9854 370574
rect 9234 334894 9854 370338
rect 9234 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 9854 334894
rect 9234 334574 9854 334658
rect 9234 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 9854 334574
rect 9234 298894 9854 334338
rect 9234 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 9854 298894
rect 9234 298574 9854 298658
rect 9234 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 9854 298574
rect 9234 262894 9854 298338
rect 9234 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 9854 262894
rect 9234 262574 9854 262658
rect 9234 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 9854 262574
rect 9234 226894 9854 262338
rect 9234 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 9854 226894
rect 9234 226574 9854 226658
rect 9234 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 9854 226574
rect 9234 190894 9854 226338
rect 9234 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 9854 190894
rect 9234 190574 9854 190658
rect 9234 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 9854 190574
rect 9234 154894 9854 190338
rect 9234 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 9854 154894
rect 9234 154574 9854 154658
rect 9234 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 9854 154574
rect 9234 118894 9854 154338
rect 9234 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 9854 118894
rect 9234 118574 9854 118658
rect 9234 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 9854 118574
rect 9234 82894 9854 118338
rect 9234 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 9854 82894
rect 9234 82574 9854 82658
rect 9234 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 9854 82574
rect 9234 46894 9854 82338
rect 9234 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 9854 46894
rect 9234 46574 9854 46658
rect 9234 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 9854 46574
rect 9234 10894 9854 46338
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect 9234 -4186 9854 10338
rect 9234 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 9854 -4186
rect 9234 -4506 9854 -4422
rect 9234 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 9854 -4506
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect 9234 -5734 9854 -4742
rect 12954 698614 13574 710042
rect 30954 711558 31574 711590
rect 30954 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 31574 711558
rect 30954 711238 31574 711322
rect 30954 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 31574 711238
rect 27234 709638 27854 709670
rect 27234 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 27854 709638
rect 27234 709318 27854 709402
rect 27234 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 27854 709318
rect 23514 707718 24134 707750
rect 23514 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 24134 707718
rect 23514 707398 24134 707482
rect 23514 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 24134 707398
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 662614 13574 698058
rect 12954 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 13574 662614
rect 12954 662294 13574 662378
rect 12954 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 13574 662294
rect 12954 626614 13574 662058
rect 12954 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 13574 626614
rect 12954 626294 13574 626378
rect 12954 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 13574 626294
rect 12954 590614 13574 626058
rect 12954 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 13574 590614
rect 12954 590294 13574 590378
rect 12954 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 13574 590294
rect 12954 554614 13574 590058
rect 12954 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 13574 554614
rect 12954 554294 13574 554378
rect 12954 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 13574 554294
rect 12954 518614 13574 554058
rect 12954 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 13574 518614
rect 12954 518294 13574 518378
rect 12954 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 13574 518294
rect 12954 482614 13574 518058
rect 12954 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 13574 482614
rect 12954 482294 13574 482378
rect 12954 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 13574 482294
rect 12954 446614 13574 482058
rect 12954 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 13574 446614
rect 12954 446294 13574 446378
rect 12954 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 13574 446294
rect 12954 410614 13574 446058
rect 12954 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 13574 410614
rect 12954 410294 13574 410378
rect 12954 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 13574 410294
rect 12954 374614 13574 410058
rect 12954 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 13574 374614
rect 12954 374294 13574 374378
rect 12954 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 13574 374294
rect 12954 338614 13574 374058
rect 12954 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 13574 338614
rect 12954 338294 13574 338378
rect 12954 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 13574 338294
rect 12954 302614 13574 338058
rect 12954 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 13574 302614
rect 12954 302294 13574 302378
rect 12954 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 13574 302294
rect 12954 266614 13574 302058
rect 12954 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 13574 266614
rect 12954 266294 13574 266378
rect 12954 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 13574 266294
rect 12954 230614 13574 266058
rect 12954 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 13574 230614
rect 12954 230294 13574 230378
rect 12954 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 13574 230294
rect 12954 194614 13574 230058
rect 12954 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 13574 194614
rect 12954 194294 13574 194378
rect 12954 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 13574 194294
rect 12954 158614 13574 194058
rect 12954 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 13574 158614
rect 12954 158294 13574 158378
rect 12954 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 13574 158294
rect 12954 122614 13574 158058
rect 12954 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 13574 122614
rect 12954 122294 13574 122378
rect 12954 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 13574 122294
rect 12954 86614 13574 122058
rect 12954 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 13574 86614
rect 12954 86294 13574 86378
rect 12954 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 13574 86294
rect 12954 50614 13574 86058
rect 12954 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 13574 50614
rect 12954 50294 13574 50378
rect 12954 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 13574 50294
rect 12954 14614 13574 50058
rect 12954 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 13574 14614
rect 12954 14294 13574 14378
rect 12954 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 13574 14294
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect 12954 -6106 13574 14058
rect 19794 705798 20414 705830
rect 19794 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 20414 705798
rect 19794 705478 20414 705562
rect 19794 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 20414 705478
rect 19794 669454 20414 705242
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -1306 20414 20898
rect 19794 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 20414 -1306
rect 19794 -1626 20414 -1542
rect 19794 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 20414 -1626
rect 19794 -1894 20414 -1862
rect 23514 673174 24134 707162
rect 23514 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 24134 673174
rect 23514 672854 24134 672938
rect 23514 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 24134 672854
rect 23514 637174 24134 672618
rect 23514 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 24134 637174
rect 23514 636854 24134 636938
rect 23514 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 24134 636854
rect 23514 601174 24134 636618
rect 23514 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 24134 601174
rect 23514 600854 24134 600938
rect 23514 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 24134 600854
rect 23514 565174 24134 600618
rect 23514 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 24134 565174
rect 23514 564854 24134 564938
rect 23514 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 24134 564854
rect 23514 529174 24134 564618
rect 23514 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 24134 529174
rect 23514 528854 24134 528938
rect 23514 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 24134 528854
rect 23514 493174 24134 528618
rect 23514 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 24134 493174
rect 23514 492854 24134 492938
rect 23514 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 24134 492854
rect 23514 457174 24134 492618
rect 23514 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 24134 457174
rect 23514 456854 24134 456938
rect 23514 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 24134 456854
rect 23514 421174 24134 456618
rect 23514 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 24134 421174
rect 23514 420854 24134 420938
rect 23514 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 24134 420854
rect 23514 385174 24134 420618
rect 23514 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 24134 385174
rect 23514 384854 24134 384938
rect 23514 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 24134 384854
rect 23514 349174 24134 384618
rect 23514 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 24134 349174
rect 23514 348854 24134 348938
rect 23514 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 24134 348854
rect 23514 313174 24134 348618
rect 23514 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 24134 313174
rect 23514 312854 24134 312938
rect 23514 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 24134 312854
rect 23514 277174 24134 312618
rect 23514 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 24134 277174
rect 23514 276854 24134 276938
rect 23514 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 24134 276854
rect 23514 241174 24134 276618
rect 23514 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 24134 241174
rect 23514 240854 24134 240938
rect 23514 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 24134 240854
rect 23514 205174 24134 240618
rect 23514 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 24134 205174
rect 23514 204854 24134 204938
rect 23514 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 24134 204854
rect 23514 169174 24134 204618
rect 23514 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 24134 169174
rect 23514 168854 24134 168938
rect 23514 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 24134 168854
rect 23514 133174 24134 168618
rect 23514 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 24134 133174
rect 23514 132854 24134 132938
rect 23514 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 24134 132854
rect 23514 97174 24134 132618
rect 23514 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 24134 97174
rect 23514 96854 24134 96938
rect 23514 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 24134 96854
rect 23514 61174 24134 96618
rect 23514 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 24134 61174
rect 23514 60854 24134 60938
rect 23514 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 24134 60854
rect 23514 25174 24134 60618
rect 23514 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 24134 25174
rect 23514 24854 24134 24938
rect 23514 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 24134 24854
rect 23514 -3226 24134 24618
rect 23514 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 24134 -3226
rect 23514 -3546 24134 -3462
rect 23514 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 24134 -3546
rect 23514 -3814 24134 -3782
rect 27234 676894 27854 709082
rect 27234 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 27854 676894
rect 27234 676574 27854 676658
rect 27234 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 27854 676574
rect 27234 640894 27854 676338
rect 27234 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 27854 640894
rect 27234 640574 27854 640658
rect 27234 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 27854 640574
rect 27234 604894 27854 640338
rect 27234 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 27854 604894
rect 27234 604574 27854 604658
rect 27234 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 27854 604574
rect 27234 568894 27854 604338
rect 27234 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 27854 568894
rect 27234 568574 27854 568658
rect 27234 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 27854 568574
rect 27234 532894 27854 568338
rect 27234 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 27854 532894
rect 27234 532574 27854 532658
rect 27234 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 27854 532574
rect 27234 496894 27854 532338
rect 27234 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 27854 496894
rect 27234 496574 27854 496658
rect 27234 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 27854 496574
rect 27234 460894 27854 496338
rect 27234 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 27854 460894
rect 27234 460574 27854 460658
rect 27234 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 27854 460574
rect 27234 424894 27854 460338
rect 27234 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 27854 424894
rect 27234 424574 27854 424658
rect 27234 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 27854 424574
rect 27234 388894 27854 424338
rect 27234 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 27854 388894
rect 27234 388574 27854 388658
rect 27234 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 27854 388574
rect 27234 352894 27854 388338
rect 27234 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 27854 352894
rect 27234 352574 27854 352658
rect 27234 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 27854 352574
rect 27234 316894 27854 352338
rect 27234 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 27854 316894
rect 27234 316574 27854 316658
rect 27234 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 27854 316574
rect 27234 280894 27854 316338
rect 27234 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 27854 280894
rect 27234 280574 27854 280658
rect 27234 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 27854 280574
rect 27234 244894 27854 280338
rect 27234 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 27854 244894
rect 27234 244574 27854 244658
rect 27234 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 27854 244574
rect 27234 208894 27854 244338
rect 27234 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 27854 208894
rect 27234 208574 27854 208658
rect 27234 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 27854 208574
rect 27234 172894 27854 208338
rect 27234 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 27854 172894
rect 27234 172574 27854 172658
rect 27234 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 27854 172574
rect 27234 136894 27854 172338
rect 27234 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 27854 136894
rect 27234 136574 27854 136658
rect 27234 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 27854 136574
rect 27234 100894 27854 136338
rect 27234 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 27854 100894
rect 27234 100574 27854 100658
rect 27234 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 27854 100574
rect 27234 64894 27854 100338
rect 27234 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 27854 64894
rect 27234 64574 27854 64658
rect 27234 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 27854 64574
rect 27234 28894 27854 64338
rect 27234 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 27854 28894
rect 27234 28574 27854 28658
rect 27234 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 27854 28574
rect 27234 -5146 27854 28338
rect 27234 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 27854 -5146
rect 27234 -5466 27854 -5382
rect 27234 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 27854 -5466
rect 27234 -5734 27854 -5702
rect 30954 680614 31574 711002
rect 48954 710598 49574 711590
rect 48954 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 49574 710598
rect 48954 710278 49574 710362
rect 48954 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 49574 710278
rect 45234 708678 45854 709670
rect 45234 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 45854 708678
rect 45234 708358 45854 708442
rect 45234 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 45854 708358
rect 41514 706758 42134 707750
rect 41514 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 42134 706758
rect 41514 706438 42134 706522
rect 41514 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 42134 706438
rect 30954 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 31574 680614
rect 30954 680294 31574 680378
rect 30954 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 31574 680294
rect 30954 644614 31574 680058
rect 30954 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 31574 644614
rect 30954 644294 31574 644378
rect 30954 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 31574 644294
rect 30954 608614 31574 644058
rect 30954 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 31574 608614
rect 30954 608294 31574 608378
rect 30954 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 31574 608294
rect 30954 572614 31574 608058
rect 30954 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 31574 572614
rect 30954 572294 31574 572378
rect 30954 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 31574 572294
rect 30954 536614 31574 572058
rect 30954 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 31574 536614
rect 30954 536294 31574 536378
rect 30954 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 31574 536294
rect 30954 500614 31574 536058
rect 30954 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 31574 500614
rect 30954 500294 31574 500378
rect 30954 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 31574 500294
rect 30954 464614 31574 500058
rect 30954 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 31574 464614
rect 30954 464294 31574 464378
rect 30954 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 31574 464294
rect 30954 428614 31574 464058
rect 30954 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 31574 428614
rect 30954 428294 31574 428378
rect 30954 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 31574 428294
rect 30954 392614 31574 428058
rect 30954 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 31574 392614
rect 30954 392294 31574 392378
rect 30954 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 31574 392294
rect 30954 356614 31574 392058
rect 30954 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 31574 356614
rect 30954 356294 31574 356378
rect 30954 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 31574 356294
rect 30954 320614 31574 356058
rect 30954 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 31574 320614
rect 30954 320294 31574 320378
rect 30954 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 31574 320294
rect 30954 284614 31574 320058
rect 30954 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 31574 284614
rect 30954 284294 31574 284378
rect 30954 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 31574 284294
rect 30954 248614 31574 284058
rect 30954 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 31574 248614
rect 30954 248294 31574 248378
rect 30954 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 31574 248294
rect 30954 212614 31574 248058
rect 30954 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 31574 212614
rect 30954 212294 31574 212378
rect 30954 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 31574 212294
rect 30954 176614 31574 212058
rect 30954 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 31574 176614
rect 30954 176294 31574 176378
rect 30954 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 31574 176294
rect 30954 140614 31574 176058
rect 30954 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 31574 140614
rect 30954 140294 31574 140378
rect 30954 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 31574 140294
rect 30954 104614 31574 140058
rect 30954 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 31574 104614
rect 30954 104294 31574 104378
rect 30954 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 31574 104294
rect 30954 68614 31574 104058
rect 30954 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 31574 68614
rect 30954 68294 31574 68378
rect 30954 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 31574 68294
rect 30954 32614 31574 68058
rect 30954 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 31574 32614
rect 30954 32294 31574 32378
rect 30954 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 31574 32294
rect 12954 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 13574 -6106
rect 12954 -6426 13574 -6342
rect 12954 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 13574 -6426
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 12954 -7654 13574 -6662
rect 30954 -7066 31574 32058
rect 37794 704838 38414 705830
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -1894 38414 -902
rect 41514 691174 42134 706202
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 41514 655174 42134 690618
rect 41514 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 42134 655174
rect 41514 654854 42134 654938
rect 41514 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 42134 654854
rect 41514 619174 42134 654618
rect 41514 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 42134 619174
rect 41514 618854 42134 618938
rect 41514 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 42134 618854
rect 41514 583174 42134 618618
rect 41514 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 42134 583174
rect 41514 582854 42134 582938
rect 41514 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 42134 582854
rect 41514 547174 42134 582618
rect 41514 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 42134 547174
rect 41514 546854 42134 546938
rect 41514 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 42134 546854
rect 41514 511174 42134 546618
rect 41514 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 42134 511174
rect 41514 510854 42134 510938
rect 41514 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 42134 510854
rect 41514 475174 42134 510618
rect 41514 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 42134 475174
rect 41514 474854 42134 474938
rect 41514 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 42134 474854
rect 41514 439174 42134 474618
rect 41514 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 42134 439174
rect 41514 438854 42134 438938
rect 41514 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 42134 438854
rect 41514 403174 42134 438618
rect 41514 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 42134 403174
rect 41514 402854 42134 402938
rect 41514 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 42134 402854
rect 41514 367174 42134 402618
rect 41514 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 42134 367174
rect 41514 366854 42134 366938
rect 41514 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 42134 366854
rect 41514 331174 42134 366618
rect 41514 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 42134 331174
rect 41514 330854 42134 330938
rect 41514 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 42134 330854
rect 41514 295174 42134 330618
rect 41514 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 42134 295174
rect 41514 294854 42134 294938
rect 41514 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 42134 294854
rect 41514 259174 42134 294618
rect 41514 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 42134 259174
rect 41514 258854 42134 258938
rect 41514 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 42134 258854
rect 41514 223174 42134 258618
rect 41514 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 42134 223174
rect 41514 222854 42134 222938
rect 41514 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 42134 222854
rect 41514 187174 42134 222618
rect 41514 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 42134 187174
rect 41514 186854 42134 186938
rect 41514 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 42134 186854
rect 41514 151174 42134 186618
rect 41514 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 42134 151174
rect 41514 150854 42134 150938
rect 41514 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 42134 150854
rect 41514 115174 42134 150618
rect 41514 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 42134 115174
rect 41514 114854 42134 114938
rect 41514 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 42134 114854
rect 41514 79174 42134 114618
rect 41514 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 42134 79174
rect 41514 78854 42134 78938
rect 41514 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 42134 78854
rect 41514 43174 42134 78618
rect 41514 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 42134 43174
rect 41514 42854 42134 42938
rect 41514 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 42134 42854
rect 41514 7174 42134 42618
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -2266 42134 6618
rect 41514 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 42134 -2266
rect 41514 -2586 42134 -2502
rect 41514 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 42134 -2586
rect 41514 -3814 42134 -2822
rect 45234 694894 45854 708122
rect 45234 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 45854 694894
rect 45234 694574 45854 694658
rect 45234 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 45854 694574
rect 45234 658894 45854 694338
rect 45234 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 45854 658894
rect 45234 658574 45854 658658
rect 45234 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 45854 658574
rect 45234 622894 45854 658338
rect 45234 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 45854 622894
rect 45234 622574 45854 622658
rect 45234 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 45854 622574
rect 45234 586894 45854 622338
rect 45234 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 45854 586894
rect 45234 586574 45854 586658
rect 45234 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 45854 586574
rect 45234 550894 45854 586338
rect 45234 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 45854 550894
rect 45234 550574 45854 550658
rect 45234 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 45854 550574
rect 45234 514894 45854 550338
rect 45234 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 45854 514894
rect 45234 514574 45854 514658
rect 45234 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 45854 514574
rect 45234 478894 45854 514338
rect 45234 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 45854 478894
rect 45234 478574 45854 478658
rect 45234 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 45854 478574
rect 45234 442894 45854 478338
rect 48954 698614 49574 710042
rect 66954 711558 67574 711590
rect 66954 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 67574 711558
rect 66954 711238 67574 711322
rect 66954 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 67574 711238
rect 63234 709638 63854 709670
rect 63234 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 63854 709638
rect 63234 709318 63854 709402
rect 63234 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 63854 709318
rect 59514 707718 60134 707750
rect 59514 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 60134 707718
rect 59514 707398 60134 707482
rect 59514 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 60134 707398
rect 48954 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 49574 698614
rect 48954 698294 49574 698378
rect 48954 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 49574 698294
rect 48954 662614 49574 698058
rect 48954 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 49574 662614
rect 48954 662294 49574 662378
rect 48954 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 49574 662294
rect 48954 626614 49574 662058
rect 48954 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 49574 626614
rect 48954 626294 49574 626378
rect 48954 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 49574 626294
rect 48954 590614 49574 626058
rect 48954 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 49574 590614
rect 48954 590294 49574 590378
rect 48954 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 49574 590294
rect 48954 554614 49574 590058
rect 48954 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 49574 554614
rect 48954 554294 49574 554378
rect 48954 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 49574 554294
rect 48954 518614 49574 554058
rect 48954 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 49574 518614
rect 48954 518294 49574 518378
rect 48954 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 49574 518294
rect 48954 482614 49574 518058
rect 48954 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 49574 482614
rect 48954 482294 49574 482378
rect 48954 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 49574 482294
rect 48954 465308 49574 482058
rect 55794 705798 56414 705830
rect 55794 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 56414 705798
rect 55794 705478 56414 705562
rect 55794 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 56414 705478
rect 55794 669454 56414 705242
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 465308 56414 488898
rect 59514 673174 60134 707162
rect 59514 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 60134 673174
rect 59514 672854 60134 672938
rect 59514 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 60134 672854
rect 59514 637174 60134 672618
rect 59514 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 60134 637174
rect 59514 636854 60134 636938
rect 59514 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 60134 636854
rect 59514 601174 60134 636618
rect 59514 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 60134 601174
rect 59514 600854 60134 600938
rect 59514 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 60134 600854
rect 59514 565174 60134 600618
rect 59514 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 60134 565174
rect 59514 564854 60134 564938
rect 59514 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 60134 564854
rect 59514 529174 60134 564618
rect 59514 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 60134 529174
rect 59514 528854 60134 528938
rect 59514 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 60134 528854
rect 59514 493174 60134 528618
rect 59514 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 60134 493174
rect 59514 492854 60134 492938
rect 59514 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 60134 492854
rect 59514 465308 60134 492618
rect 63234 676894 63854 709082
rect 63234 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 63854 676894
rect 63234 676574 63854 676658
rect 63234 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 63854 676574
rect 63234 640894 63854 676338
rect 63234 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 63854 640894
rect 63234 640574 63854 640658
rect 63234 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 63854 640574
rect 63234 604894 63854 640338
rect 63234 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 63854 604894
rect 63234 604574 63854 604658
rect 63234 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 63854 604574
rect 63234 568894 63854 604338
rect 63234 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 63854 568894
rect 63234 568574 63854 568658
rect 63234 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 63854 568574
rect 63234 532894 63854 568338
rect 63234 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 63854 532894
rect 63234 532574 63854 532658
rect 63234 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 63854 532574
rect 63234 496894 63854 532338
rect 63234 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 63854 496894
rect 63234 496574 63854 496658
rect 63234 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 63854 496574
rect 63234 465308 63854 496338
rect 66954 680614 67574 711002
rect 84954 710598 85574 711590
rect 84954 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 85574 710598
rect 84954 710278 85574 710362
rect 84954 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 85574 710278
rect 81234 708678 81854 709670
rect 81234 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 81854 708678
rect 81234 708358 81854 708442
rect 81234 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 81854 708358
rect 77514 706758 78134 707750
rect 77514 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 78134 706758
rect 77514 706438 78134 706522
rect 77514 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 78134 706438
rect 66954 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 67574 680614
rect 66954 680294 67574 680378
rect 66954 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 67574 680294
rect 66954 644614 67574 680058
rect 66954 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 67574 644614
rect 66954 644294 67574 644378
rect 66954 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 67574 644294
rect 66954 608614 67574 644058
rect 66954 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 67574 608614
rect 66954 608294 67574 608378
rect 66954 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 67574 608294
rect 66954 572614 67574 608058
rect 66954 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 67574 572614
rect 66954 572294 67574 572378
rect 66954 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 67574 572294
rect 66954 536614 67574 572058
rect 66954 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 67574 536614
rect 66954 536294 67574 536378
rect 66954 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 67574 536294
rect 66954 500614 67574 536058
rect 66954 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 67574 500614
rect 66954 500294 67574 500378
rect 66954 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 67574 500294
rect 66954 465308 67574 500058
rect 73794 704838 74414 705830
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 579454 74414 614898
rect 73794 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 74414 579454
rect 73794 579134 74414 579218
rect 73794 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 74414 579134
rect 73794 543454 74414 578898
rect 73794 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 74414 543454
rect 73794 543134 74414 543218
rect 73794 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 74414 543134
rect 73794 507454 74414 542898
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 471454 74414 506898
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73794 465308 74414 470898
rect 77514 691174 78134 706202
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 655174 78134 690618
rect 77514 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 78134 655174
rect 77514 654854 78134 654938
rect 77514 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 78134 654854
rect 77514 619174 78134 654618
rect 77514 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 78134 619174
rect 77514 618854 78134 618938
rect 77514 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 78134 618854
rect 77514 583174 78134 618618
rect 77514 582938 77546 583174
rect 77782 582938 77866 583174
rect 78102 582938 78134 583174
rect 77514 582854 78134 582938
rect 77514 582618 77546 582854
rect 77782 582618 77866 582854
rect 78102 582618 78134 582854
rect 77514 547174 78134 582618
rect 77514 546938 77546 547174
rect 77782 546938 77866 547174
rect 78102 546938 78134 547174
rect 77514 546854 78134 546938
rect 77514 546618 77546 546854
rect 77782 546618 77866 546854
rect 78102 546618 78134 546854
rect 77514 511174 78134 546618
rect 77514 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 78134 511174
rect 77514 510854 78134 510938
rect 77514 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 78134 510854
rect 77514 475174 78134 510618
rect 77514 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 78134 475174
rect 77514 474854 78134 474938
rect 77514 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 78134 474854
rect 77514 465308 78134 474618
rect 81234 694894 81854 708122
rect 81234 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 81854 694894
rect 81234 694574 81854 694658
rect 81234 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 81854 694574
rect 81234 658894 81854 694338
rect 81234 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 81854 658894
rect 81234 658574 81854 658658
rect 81234 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 81854 658574
rect 81234 622894 81854 658338
rect 81234 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 81854 622894
rect 81234 622574 81854 622658
rect 81234 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 81854 622574
rect 81234 586894 81854 622338
rect 81234 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 81854 586894
rect 81234 586574 81854 586658
rect 81234 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 81854 586574
rect 81234 550894 81854 586338
rect 81234 550658 81266 550894
rect 81502 550658 81586 550894
rect 81822 550658 81854 550894
rect 81234 550574 81854 550658
rect 81234 550338 81266 550574
rect 81502 550338 81586 550574
rect 81822 550338 81854 550574
rect 81234 514894 81854 550338
rect 81234 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 81854 514894
rect 81234 514574 81854 514658
rect 81234 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 81854 514574
rect 81234 478894 81854 514338
rect 81234 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 81854 478894
rect 81234 478574 81854 478658
rect 81234 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 81854 478574
rect 81019 465628 81085 465629
rect 81019 465564 81020 465628
rect 81084 465564 81085 465628
rect 81019 465563 81085 465564
rect 78811 465356 78877 465357
rect 78811 465292 78812 465356
rect 78876 465292 78877 465356
rect 78811 465291 78877 465292
rect 78814 463450 78874 465291
rect 81022 463450 81082 465563
rect 81234 465308 81854 478338
rect 84954 698614 85574 710042
rect 102954 711558 103574 711590
rect 102954 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 103574 711558
rect 102954 711238 103574 711322
rect 102954 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 103574 711238
rect 99234 709638 99854 709670
rect 99234 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 99854 709638
rect 99234 709318 99854 709402
rect 99234 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 99854 709318
rect 95514 707718 96134 707750
rect 95514 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 96134 707718
rect 95514 707398 96134 707482
rect 95514 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 96134 707398
rect 84954 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 85574 698614
rect 84954 698294 85574 698378
rect 84954 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 85574 698294
rect 84954 662614 85574 698058
rect 84954 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 85574 662614
rect 84954 662294 85574 662378
rect 84954 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 85574 662294
rect 84954 626614 85574 662058
rect 84954 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 85574 626614
rect 84954 626294 85574 626378
rect 84954 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 85574 626294
rect 84954 590614 85574 626058
rect 84954 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 85574 590614
rect 84954 590294 85574 590378
rect 84954 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 85574 590294
rect 84954 554614 85574 590058
rect 84954 554378 84986 554614
rect 85222 554378 85306 554614
rect 85542 554378 85574 554614
rect 84954 554294 85574 554378
rect 84954 554058 84986 554294
rect 85222 554058 85306 554294
rect 85542 554058 85574 554294
rect 84954 518614 85574 554058
rect 84954 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 85574 518614
rect 84954 518294 85574 518378
rect 84954 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 85574 518294
rect 84954 482614 85574 518058
rect 84954 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 85574 482614
rect 84954 482294 85574 482378
rect 84954 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 85574 482294
rect 84954 465308 85574 482058
rect 91794 705798 92414 705830
rect 91794 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 92414 705798
rect 91794 705478 92414 705562
rect 91794 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 92414 705478
rect 91794 669454 92414 705242
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 91794 561454 92414 596898
rect 91794 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 92414 561454
rect 91794 561134 92414 561218
rect 91794 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 92414 561134
rect 91794 525454 92414 560898
rect 91794 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 92414 525454
rect 91794 525134 92414 525218
rect 91794 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 92414 525134
rect 91794 489454 92414 524898
rect 91794 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 92414 489454
rect 91794 489134 92414 489218
rect 91794 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 92414 489134
rect 86171 465492 86237 465493
rect 86171 465428 86172 465492
rect 86236 465428 86237 465492
rect 86171 465427 86237 465428
rect 83461 463724 83527 463725
rect 83461 463660 83462 463724
rect 83526 463660 83527 463724
rect 83461 463659 83527 463660
rect 78704 463390 78874 463450
rect 81016 463390 81082 463450
rect 78704 463202 78764 463390
rect 81016 463202 81076 463390
rect 83464 463202 83524 463659
rect 86174 463450 86234 465427
rect 91794 465308 92414 488898
rect 95514 673174 96134 707162
rect 95514 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 96134 673174
rect 95514 672854 96134 672938
rect 95514 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 96134 672854
rect 95514 637174 96134 672618
rect 95514 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 96134 637174
rect 95514 636854 96134 636938
rect 95514 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 96134 636854
rect 95514 601174 96134 636618
rect 95514 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 96134 601174
rect 95514 600854 96134 600938
rect 95514 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 96134 600854
rect 95514 565174 96134 600618
rect 95514 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 96134 565174
rect 95514 564854 96134 564938
rect 95514 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 96134 564854
rect 95514 529174 96134 564618
rect 95514 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 96134 529174
rect 95514 528854 96134 528938
rect 95514 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 96134 528854
rect 95514 493174 96134 528618
rect 95514 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 96134 493174
rect 95514 492854 96134 492938
rect 95514 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 96134 492854
rect 95514 465308 96134 492618
rect 99234 676894 99854 709082
rect 99234 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 99854 676894
rect 99234 676574 99854 676658
rect 99234 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 99854 676574
rect 99234 640894 99854 676338
rect 99234 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 99854 640894
rect 99234 640574 99854 640658
rect 99234 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 99854 640574
rect 99234 604894 99854 640338
rect 99234 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 99854 604894
rect 99234 604574 99854 604658
rect 99234 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 99854 604574
rect 99234 568894 99854 604338
rect 99234 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 99854 568894
rect 99234 568574 99854 568658
rect 99234 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 99854 568574
rect 99234 532894 99854 568338
rect 99234 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 99854 532894
rect 99234 532574 99854 532658
rect 99234 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 99854 532574
rect 99234 496894 99854 532338
rect 99234 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 99854 496894
rect 99234 496574 99854 496658
rect 99234 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 99854 496574
rect 99234 465308 99854 496338
rect 102954 680614 103574 711002
rect 120954 710598 121574 711590
rect 120954 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 121574 710598
rect 120954 710278 121574 710362
rect 120954 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 121574 710278
rect 117234 708678 117854 709670
rect 117234 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 117854 708678
rect 117234 708358 117854 708442
rect 117234 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 117854 708358
rect 113514 706758 114134 707750
rect 113514 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 114134 706758
rect 113514 706438 114134 706522
rect 113514 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 114134 706438
rect 102954 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 103574 680614
rect 102954 680294 103574 680378
rect 102954 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 103574 680294
rect 102954 644614 103574 680058
rect 102954 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 103574 644614
rect 102954 644294 103574 644378
rect 102954 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 103574 644294
rect 102954 608614 103574 644058
rect 102954 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 103574 608614
rect 102954 608294 103574 608378
rect 102954 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 103574 608294
rect 102954 572614 103574 608058
rect 102954 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 103574 572614
rect 102954 572294 103574 572378
rect 102954 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 103574 572294
rect 102954 536614 103574 572058
rect 102954 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 103574 536614
rect 102954 536294 103574 536378
rect 102954 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 103574 536294
rect 102954 500614 103574 536058
rect 102954 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 103574 500614
rect 102954 500294 103574 500378
rect 102954 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 103574 500294
rect 102954 465308 103574 500058
rect 109794 704838 110414 705830
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 109794 543454 110414 578898
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 109794 507454 110414 542898
rect 109794 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 110414 507454
rect 109794 507134 110414 507218
rect 109794 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 110414 507134
rect 109794 471454 110414 506898
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 109794 465308 110414 470898
rect 113514 691174 114134 706202
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 113514 655174 114134 690618
rect 113514 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 114134 655174
rect 113514 654854 114134 654938
rect 113514 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 114134 654854
rect 113514 619174 114134 654618
rect 113514 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 114134 619174
rect 113514 618854 114134 618938
rect 113514 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 114134 618854
rect 113514 583174 114134 618618
rect 113514 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 114134 583174
rect 113514 582854 114134 582938
rect 113514 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 114134 582854
rect 113514 547174 114134 582618
rect 113514 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 114134 547174
rect 113514 546854 114134 546938
rect 113514 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 114134 546854
rect 113514 511174 114134 546618
rect 113514 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 114134 511174
rect 113514 510854 114134 510938
rect 113514 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 114134 510854
rect 113514 475174 114134 510618
rect 113514 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 114134 475174
rect 113514 474854 114134 474938
rect 113514 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 114134 474854
rect 113514 465308 114134 474618
rect 117234 694894 117854 708122
rect 117234 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 117854 694894
rect 117234 694574 117854 694658
rect 117234 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 117854 694574
rect 117234 658894 117854 694338
rect 117234 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 117854 658894
rect 117234 658574 117854 658658
rect 117234 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 117854 658574
rect 117234 622894 117854 658338
rect 117234 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 117854 622894
rect 117234 622574 117854 622658
rect 117234 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 117854 622574
rect 117234 586894 117854 622338
rect 117234 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 117854 586894
rect 117234 586574 117854 586658
rect 117234 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 117854 586574
rect 117234 550894 117854 586338
rect 117234 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 117854 550894
rect 117234 550574 117854 550658
rect 117234 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 117854 550574
rect 117234 514894 117854 550338
rect 117234 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 117854 514894
rect 117234 514574 117854 514658
rect 117234 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 117854 514574
rect 117234 478894 117854 514338
rect 117234 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 117854 478894
rect 117234 478574 117854 478658
rect 117234 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 117854 478574
rect 117234 465308 117854 478338
rect 120954 698614 121574 710042
rect 138954 711558 139574 711590
rect 138954 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 139574 711558
rect 138954 711238 139574 711322
rect 138954 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 139574 711238
rect 135234 709638 135854 709670
rect 135234 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 135854 709638
rect 135234 709318 135854 709402
rect 135234 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 135854 709318
rect 131514 707718 132134 707750
rect 131514 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 132134 707718
rect 131514 707398 132134 707482
rect 131514 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 132134 707398
rect 120954 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 121574 698614
rect 120954 698294 121574 698378
rect 120954 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 121574 698294
rect 120954 662614 121574 698058
rect 120954 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 121574 662614
rect 120954 662294 121574 662378
rect 120954 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 121574 662294
rect 120954 626614 121574 662058
rect 120954 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 121574 626614
rect 120954 626294 121574 626378
rect 120954 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 121574 626294
rect 120954 590614 121574 626058
rect 120954 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 121574 590614
rect 120954 590294 121574 590378
rect 120954 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 121574 590294
rect 120954 554614 121574 590058
rect 120954 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 121574 554614
rect 120954 554294 121574 554378
rect 120954 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 121574 554294
rect 120954 518614 121574 554058
rect 120954 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 121574 518614
rect 120954 518294 121574 518378
rect 120954 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 121574 518294
rect 120954 482614 121574 518058
rect 120954 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 121574 482614
rect 120954 482294 121574 482378
rect 120954 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 121574 482294
rect 120954 465308 121574 482058
rect 127794 705798 128414 705830
rect 127794 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 128414 705798
rect 127794 705478 128414 705562
rect 127794 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 128414 705478
rect 127794 669454 128414 705242
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 127794 561454 128414 596898
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 127794 525454 128414 560898
rect 127794 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 128414 525454
rect 127794 525134 128414 525218
rect 127794 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 128414 525134
rect 127794 489454 128414 524898
rect 127794 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 128414 489454
rect 127794 489134 128414 489218
rect 127794 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 128414 489134
rect 127794 465308 128414 488898
rect 131514 673174 132134 707162
rect 131514 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 132134 673174
rect 131514 672854 132134 672938
rect 131514 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 132134 672854
rect 131514 637174 132134 672618
rect 131514 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 132134 637174
rect 131514 636854 132134 636938
rect 131514 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 132134 636854
rect 131514 601174 132134 636618
rect 131514 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 132134 601174
rect 131514 600854 132134 600938
rect 131514 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 132134 600854
rect 131514 565174 132134 600618
rect 131514 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 132134 565174
rect 131514 564854 132134 564938
rect 131514 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 132134 564854
rect 131514 529174 132134 564618
rect 131514 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 132134 529174
rect 131514 528854 132134 528938
rect 131514 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 132134 528854
rect 131514 493174 132134 528618
rect 131514 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 132134 493174
rect 131514 492854 132134 492938
rect 131514 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 132134 492854
rect 131514 465308 132134 492618
rect 135234 676894 135854 709082
rect 135234 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 135854 676894
rect 135234 676574 135854 676658
rect 135234 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 135854 676574
rect 135234 640894 135854 676338
rect 135234 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 135854 640894
rect 135234 640574 135854 640658
rect 135234 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 135854 640574
rect 135234 604894 135854 640338
rect 135234 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 135854 604894
rect 135234 604574 135854 604658
rect 135234 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 135854 604574
rect 135234 568894 135854 604338
rect 135234 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 135854 568894
rect 135234 568574 135854 568658
rect 135234 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 135854 568574
rect 135234 532894 135854 568338
rect 135234 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 135854 532894
rect 135234 532574 135854 532658
rect 135234 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 135854 532574
rect 135234 496894 135854 532338
rect 135234 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 135854 496894
rect 135234 496574 135854 496658
rect 135234 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 135854 496574
rect 135234 465308 135854 496338
rect 138954 680614 139574 711002
rect 156954 710598 157574 711590
rect 156954 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 157574 710598
rect 156954 710278 157574 710362
rect 156954 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 157574 710278
rect 153234 708678 153854 709670
rect 153234 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 153854 708678
rect 153234 708358 153854 708442
rect 153234 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 153854 708358
rect 149514 706758 150134 707750
rect 149514 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 150134 706758
rect 149514 706438 150134 706522
rect 149514 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 150134 706438
rect 138954 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 139574 680614
rect 138954 680294 139574 680378
rect 138954 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 139574 680294
rect 138954 644614 139574 680058
rect 138954 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 139574 644614
rect 138954 644294 139574 644378
rect 138954 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 139574 644294
rect 138954 608614 139574 644058
rect 138954 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 139574 608614
rect 138954 608294 139574 608378
rect 138954 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 139574 608294
rect 138954 572614 139574 608058
rect 138954 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 139574 572614
rect 138954 572294 139574 572378
rect 138954 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 139574 572294
rect 138954 536614 139574 572058
rect 138954 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 139574 536614
rect 138954 536294 139574 536378
rect 138954 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 139574 536294
rect 138954 500614 139574 536058
rect 138954 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 139574 500614
rect 138954 500294 139574 500378
rect 138954 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 139574 500294
rect 138954 465308 139574 500058
rect 145794 704838 146414 705830
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 543454 146414 578898
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 507454 146414 542898
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 145794 471454 146414 506898
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 465308 146414 470898
rect 149514 691174 150134 706202
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 655174 150134 690618
rect 149514 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 150134 655174
rect 149514 654854 150134 654938
rect 149514 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 150134 654854
rect 149514 619174 150134 654618
rect 149514 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 150134 619174
rect 149514 618854 150134 618938
rect 149514 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 150134 618854
rect 149514 583174 150134 618618
rect 149514 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 150134 583174
rect 149514 582854 150134 582938
rect 149514 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 150134 582854
rect 149514 547174 150134 582618
rect 149514 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 150134 547174
rect 149514 546854 150134 546938
rect 149514 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 150134 546854
rect 149514 511174 150134 546618
rect 149514 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 150134 511174
rect 149514 510854 150134 510938
rect 149514 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 150134 510854
rect 149514 475174 150134 510618
rect 149514 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 150134 475174
rect 149514 474854 150134 474938
rect 149514 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 150134 474854
rect 149514 465308 150134 474618
rect 153234 694894 153854 708122
rect 153234 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 153854 694894
rect 153234 694574 153854 694658
rect 153234 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 153854 694574
rect 153234 658894 153854 694338
rect 153234 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 153854 658894
rect 153234 658574 153854 658658
rect 153234 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 153854 658574
rect 153234 622894 153854 658338
rect 153234 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 153854 622894
rect 153234 622574 153854 622658
rect 153234 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 153854 622574
rect 153234 586894 153854 622338
rect 153234 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 153854 586894
rect 153234 586574 153854 586658
rect 153234 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 153854 586574
rect 153234 550894 153854 586338
rect 153234 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 153854 550894
rect 153234 550574 153854 550658
rect 153234 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 153854 550574
rect 153234 514894 153854 550338
rect 153234 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 153854 514894
rect 153234 514574 153854 514658
rect 153234 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 153854 514574
rect 153234 478894 153854 514338
rect 153234 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 153854 478894
rect 153234 478574 153854 478658
rect 153234 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 153854 478574
rect 151123 466308 151189 466309
rect 151123 466244 151124 466308
rect 151188 466244 151189 466308
rect 151123 466243 151189 466244
rect 91139 465220 91205 465221
rect 91139 465156 91140 465220
rect 91204 465156 91205 465220
rect 91139 465155 91205 465156
rect 93531 465220 93597 465221
rect 93531 465156 93532 465220
rect 93596 465156 93597 465220
rect 93531 465155 93597 465156
rect 96107 465220 96173 465221
rect 96107 465156 96108 465220
rect 96172 465156 96173 465220
rect 96107 465155 96173 465156
rect 101259 465220 101325 465221
rect 101259 465156 101260 465220
rect 101324 465156 101325 465220
rect 101259 465155 101325 465156
rect 103651 465220 103717 465221
rect 103651 465156 103652 465220
rect 103716 465156 103717 465220
rect 103651 465155 103717 465156
rect 106227 465220 106293 465221
rect 106227 465156 106228 465220
rect 106292 465156 106293 465220
rect 106227 465155 106293 465156
rect 108435 465220 108501 465221
rect 108435 465156 108436 465220
rect 108500 465156 108501 465220
rect 108435 465155 108501 465156
rect 111011 465220 111077 465221
rect 111011 465156 111012 465220
rect 111076 465156 111077 465220
rect 111011 465155 111077 465156
rect 128675 465220 128741 465221
rect 128675 465156 128676 465220
rect 128740 465156 128741 465220
rect 128675 465155 128741 465156
rect 136035 465220 136101 465221
rect 136035 465156 136036 465220
rect 136100 465156 136101 465220
rect 136035 465155 136101 465156
rect 141003 465220 141069 465221
rect 141003 465156 141004 465220
rect 141068 465156 141069 465220
rect 141003 465155 141069 465156
rect 145971 465220 146037 465221
rect 145971 465156 145972 465220
rect 146036 465156 146037 465220
rect 145971 465155 146037 465156
rect 88493 463724 88559 463725
rect 88493 463660 88494 463724
rect 88558 463660 88559 463724
rect 88493 463659 88559 463660
rect 86174 463390 86244 463450
rect 86184 463202 86244 463390
rect 88496 463202 88556 463659
rect 91142 463450 91202 465155
rect 93534 463450 93594 465155
rect 96110 463710 96170 465155
rect 98557 463724 98623 463725
rect 96110 463650 96172 463710
rect 98557 463660 98558 463724
rect 98622 463660 98623 463724
rect 101262 463710 101322 465155
rect 98557 463659 98623 463660
rect 91080 463390 91202 463450
rect 93528 463390 93594 463450
rect 91080 463202 91140 463390
rect 93528 463202 93588 463390
rect 96112 463202 96172 463650
rect 98560 463202 98620 463659
rect 101144 463650 101322 463710
rect 101144 463202 101204 463650
rect 103654 463450 103714 465155
rect 106230 463450 106290 465155
rect 103592 463390 103714 463450
rect 106176 463390 106290 463450
rect 108438 463450 108498 465155
rect 111014 463450 111074 465155
rect 113653 463724 113719 463725
rect 113653 463660 113654 463724
rect 113718 463660 113719 463724
rect 113653 463659 113719 463660
rect 116101 463724 116167 463725
rect 116101 463660 116102 463724
rect 116166 463660 116167 463724
rect 116101 463659 116167 463660
rect 118549 463724 118615 463725
rect 118549 463660 118550 463724
rect 118614 463660 118615 463724
rect 118549 463659 118615 463660
rect 120997 463724 121063 463725
rect 120997 463660 120998 463724
rect 121062 463660 121063 463724
rect 120997 463659 121063 463660
rect 123581 463724 123647 463725
rect 123581 463660 123582 463724
rect 123646 463660 123647 463724
rect 123581 463659 123647 463660
rect 125893 463724 125959 463725
rect 125893 463660 125894 463724
rect 125958 463660 125959 463724
rect 125893 463659 125959 463660
rect 108438 463390 108548 463450
rect 103592 463202 103652 463390
rect 106176 463202 106236 463390
rect 108488 463202 108548 463390
rect 110936 463390 111074 463450
rect 110936 463202 110996 463390
rect 113656 463202 113716 463659
rect 116104 463202 116164 463659
rect 118552 463202 118612 463659
rect 121000 463202 121060 463659
rect 123584 463202 123644 463659
rect 125896 463202 125956 463659
rect 128678 463450 128738 465155
rect 131067 463996 131133 463997
rect 131067 463932 131068 463996
rect 131132 463932 131133 463996
rect 131067 463931 131133 463932
rect 131070 463450 131130 463931
rect 133509 463724 133575 463725
rect 133509 463660 133510 463724
rect 133574 463660 133575 463724
rect 133509 463659 133575 463660
rect 128616 463390 128738 463450
rect 131064 463390 131130 463450
rect 128616 463202 128676 463390
rect 131064 463202 131124 463390
rect 133512 463202 133572 463659
rect 136038 463450 136098 465155
rect 138405 463724 138471 463725
rect 138405 463660 138406 463724
rect 138470 463660 138471 463724
rect 138405 463659 138471 463660
rect 135960 463390 136098 463450
rect 135960 463202 136020 463390
rect 138408 463202 138468 463659
rect 141006 463450 141066 465155
rect 143573 463724 143639 463725
rect 143573 463660 143574 463724
rect 143638 463660 143639 463724
rect 143573 463659 143639 463660
rect 140992 463390 141066 463450
rect 140992 463202 141052 463390
rect 143576 463202 143636 463659
rect 145974 463450 146034 465155
rect 148469 463724 148535 463725
rect 148469 463660 148470 463724
rect 148534 463660 148535 463724
rect 148469 463659 148535 463660
rect 145974 463390 146084 463450
rect 146024 463202 146084 463390
rect 148472 463202 148532 463659
rect 151126 463450 151186 466243
rect 153234 465308 153854 478338
rect 156954 698614 157574 710042
rect 174954 711558 175574 711590
rect 174954 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 175574 711558
rect 174954 711238 175574 711322
rect 174954 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 175574 711238
rect 171234 709638 171854 709670
rect 171234 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 171854 709638
rect 171234 709318 171854 709402
rect 171234 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 171854 709318
rect 167514 707718 168134 707750
rect 167514 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 168134 707718
rect 167514 707398 168134 707482
rect 167514 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 168134 707398
rect 156954 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 157574 698614
rect 156954 698294 157574 698378
rect 156954 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 157574 698294
rect 156954 662614 157574 698058
rect 156954 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 157574 662614
rect 156954 662294 157574 662378
rect 156954 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 157574 662294
rect 156954 626614 157574 662058
rect 156954 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 157574 626614
rect 156954 626294 157574 626378
rect 156954 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 157574 626294
rect 156954 590614 157574 626058
rect 156954 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 157574 590614
rect 156954 590294 157574 590378
rect 156954 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 157574 590294
rect 156954 554614 157574 590058
rect 156954 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 157574 554614
rect 156954 554294 157574 554378
rect 156954 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 157574 554294
rect 156954 518614 157574 554058
rect 156954 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 157574 518614
rect 156954 518294 157574 518378
rect 156954 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 157574 518294
rect 156954 482614 157574 518058
rect 156954 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 157574 482614
rect 156954 482294 157574 482378
rect 156954 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 157574 482294
rect 156091 466444 156157 466445
rect 156091 466380 156092 466444
rect 156156 466380 156157 466444
rect 156091 466379 156157 466380
rect 153331 465220 153397 465221
rect 153331 465156 153332 465220
rect 153396 465156 153397 465220
rect 153331 465155 153397 465156
rect 151056 463390 151186 463450
rect 153334 463450 153394 465155
rect 156094 463450 156154 466379
rect 156954 465308 157574 482058
rect 163794 705798 164414 705830
rect 163794 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 164414 705798
rect 163794 705478 164414 705562
rect 163794 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 164414 705478
rect 163794 669454 164414 705242
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 163794 561454 164414 596898
rect 163794 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 164414 561454
rect 163794 561134 164414 561218
rect 163794 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 164414 561134
rect 163794 525454 164414 560898
rect 163794 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 164414 525454
rect 163794 525134 164414 525218
rect 163794 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 164414 525134
rect 163794 489454 164414 524898
rect 163794 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 164414 489454
rect 163794 489134 164414 489218
rect 163794 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 164414 489134
rect 163794 465308 164414 488898
rect 167514 673174 168134 707162
rect 167514 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 168134 673174
rect 167514 672854 168134 672938
rect 167514 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 168134 672854
rect 167514 637174 168134 672618
rect 167514 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 168134 637174
rect 167514 636854 168134 636938
rect 167514 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 168134 636854
rect 167514 601174 168134 636618
rect 167514 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 168134 601174
rect 167514 600854 168134 600938
rect 167514 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 168134 600854
rect 167514 565174 168134 600618
rect 167514 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 168134 565174
rect 167514 564854 168134 564938
rect 167514 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 168134 564854
rect 167514 529174 168134 564618
rect 167514 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 168134 529174
rect 167514 528854 168134 528938
rect 167514 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 168134 528854
rect 167514 493174 168134 528618
rect 167514 492938 167546 493174
rect 167782 492938 167866 493174
rect 168102 492938 168134 493174
rect 167514 492854 168134 492938
rect 167514 492618 167546 492854
rect 167782 492618 167866 492854
rect 168102 492618 168134 492854
rect 167514 465308 168134 492618
rect 171234 676894 171854 709082
rect 171234 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 171854 676894
rect 171234 676574 171854 676658
rect 171234 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 171854 676574
rect 171234 640894 171854 676338
rect 171234 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 171854 640894
rect 171234 640574 171854 640658
rect 171234 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 171854 640574
rect 171234 604894 171854 640338
rect 171234 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 171854 604894
rect 171234 604574 171854 604658
rect 171234 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 171854 604574
rect 171234 568894 171854 604338
rect 171234 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 171854 568894
rect 171234 568574 171854 568658
rect 171234 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 171854 568574
rect 171234 532894 171854 568338
rect 171234 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 171854 532894
rect 171234 532574 171854 532658
rect 171234 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 171854 532574
rect 171234 496894 171854 532338
rect 171234 496658 171266 496894
rect 171502 496658 171586 496894
rect 171822 496658 171854 496894
rect 171234 496574 171854 496658
rect 171234 496338 171266 496574
rect 171502 496338 171586 496574
rect 171822 496338 171854 496574
rect 171234 465308 171854 496338
rect 174954 680614 175574 711002
rect 192954 710598 193574 711590
rect 192954 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 193574 710598
rect 192954 710278 193574 710362
rect 192954 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 193574 710278
rect 189234 708678 189854 709670
rect 189234 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 189854 708678
rect 189234 708358 189854 708442
rect 189234 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 189854 708358
rect 185514 706758 186134 707750
rect 185514 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 186134 706758
rect 185514 706438 186134 706522
rect 185514 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 186134 706438
rect 174954 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 175574 680614
rect 174954 680294 175574 680378
rect 174954 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 175574 680294
rect 174954 644614 175574 680058
rect 174954 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 175574 644614
rect 174954 644294 175574 644378
rect 174954 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 175574 644294
rect 174954 608614 175574 644058
rect 174954 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 175574 608614
rect 174954 608294 175574 608378
rect 174954 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 175574 608294
rect 174954 572614 175574 608058
rect 174954 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 175574 572614
rect 174954 572294 175574 572378
rect 174954 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 175574 572294
rect 174954 536614 175574 572058
rect 174954 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 175574 536614
rect 174954 536294 175574 536378
rect 174954 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 175574 536294
rect 174954 500614 175574 536058
rect 174954 500378 174986 500614
rect 175222 500378 175306 500614
rect 175542 500378 175574 500614
rect 174954 500294 175574 500378
rect 174954 500058 174986 500294
rect 175222 500058 175306 500294
rect 175542 500058 175574 500294
rect 174954 465308 175574 500058
rect 181794 704838 182414 705830
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 181794 471454 182414 506898
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 181794 465308 182414 470898
rect 185514 691174 186134 706202
rect 185514 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 186134 691174
rect 185514 690854 186134 690938
rect 185514 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 186134 690854
rect 185514 655174 186134 690618
rect 185514 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 186134 655174
rect 185514 654854 186134 654938
rect 185514 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 186134 654854
rect 185514 619174 186134 654618
rect 185514 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 186134 619174
rect 185514 618854 186134 618938
rect 185514 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 186134 618854
rect 185514 583174 186134 618618
rect 185514 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 186134 583174
rect 185514 582854 186134 582938
rect 185514 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 186134 582854
rect 185514 547174 186134 582618
rect 185514 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 186134 547174
rect 185514 546854 186134 546938
rect 185514 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 186134 546854
rect 185514 511174 186134 546618
rect 185514 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 186134 511174
rect 185514 510854 186134 510938
rect 185514 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 186134 510854
rect 185514 475174 186134 510618
rect 185514 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 186134 475174
rect 185514 474854 186134 474938
rect 185514 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 186134 474854
rect 185514 465308 186134 474618
rect 189234 694894 189854 708122
rect 189234 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 189854 694894
rect 189234 694574 189854 694658
rect 189234 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 189854 694574
rect 189234 658894 189854 694338
rect 189234 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 189854 658894
rect 189234 658574 189854 658658
rect 189234 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 189854 658574
rect 189234 622894 189854 658338
rect 189234 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 189854 622894
rect 189234 622574 189854 622658
rect 189234 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 189854 622574
rect 189234 586894 189854 622338
rect 189234 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 189854 586894
rect 189234 586574 189854 586658
rect 189234 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 189854 586574
rect 189234 550894 189854 586338
rect 189234 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 189854 550894
rect 189234 550574 189854 550658
rect 189234 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 189854 550574
rect 189234 514894 189854 550338
rect 189234 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 189854 514894
rect 189234 514574 189854 514658
rect 189234 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 189854 514574
rect 189234 478894 189854 514338
rect 189234 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 189854 478894
rect 189234 478574 189854 478658
rect 189234 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 189854 478574
rect 188291 465356 188357 465357
rect 188291 465292 188292 465356
rect 188356 465292 188357 465356
rect 188291 465291 188357 465292
rect 168419 465220 168485 465221
rect 168419 465156 168420 465220
rect 168484 465156 168485 465220
rect 168419 465155 168485 465156
rect 169707 465220 169773 465221
rect 169707 465156 169708 465220
rect 169772 465156 169773 465220
rect 169707 465155 169773 465156
rect 180931 465220 180997 465221
rect 180931 465156 180932 465220
rect 180996 465156 180997 465220
rect 180931 465155 180997 465156
rect 187739 465220 187805 465221
rect 187739 465156 187740 465220
rect 187804 465156 187805 465220
rect 187739 465155 187805 465156
rect 153334 463390 153428 463450
rect 151056 463202 151116 463390
rect 153368 463202 153428 463390
rect 156088 463390 156154 463450
rect 168422 463450 168482 465155
rect 169710 463450 169770 465155
rect 180934 463450 180994 465155
rect 168422 463390 168524 463450
rect 156088 463202 156148 463390
rect 168464 463202 168524 463390
rect 169688 463390 169770 463450
rect 180840 463390 180994 463450
rect 169688 463202 169748 463390
rect 180840 463202 180900 463390
rect 186819 461004 186885 461005
rect 186819 460940 186820 461004
rect 186884 460940 186885 461004
rect 186819 460939 186885 460940
rect 50272 453454 50620 453486
rect 50272 453218 50328 453454
rect 50564 453218 50620 453454
rect 50272 453134 50620 453218
rect 50272 452898 50328 453134
rect 50564 452898 50620 453134
rect 50272 452866 50620 452898
rect 186000 453454 186348 453486
rect 186000 453218 186056 453454
rect 186292 453218 186348 453454
rect 186000 453134 186348 453218
rect 186000 452898 186056 453134
rect 186292 452898 186348 453134
rect 186000 452866 186348 452898
rect 45234 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 45854 442894
rect 45234 442574 45854 442658
rect 45234 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 45854 442574
rect 45234 406894 45854 442338
rect 50952 435454 51300 435486
rect 50952 435218 51008 435454
rect 51244 435218 51300 435454
rect 50952 435134 51300 435218
rect 50952 434898 51008 435134
rect 51244 434898 51300 435134
rect 50952 434866 51300 434898
rect 185320 435454 185668 435486
rect 185320 435218 185376 435454
rect 185612 435218 185668 435454
rect 185320 435134 185668 435218
rect 185320 434898 185376 435134
rect 185612 434898 185668 435134
rect 185320 434866 185668 434898
rect 50272 417454 50620 417486
rect 50272 417218 50328 417454
rect 50564 417218 50620 417454
rect 50272 417134 50620 417218
rect 50272 416898 50328 417134
rect 50564 416898 50620 417134
rect 50272 416866 50620 416898
rect 186000 417454 186348 417486
rect 186000 417218 186056 417454
rect 186292 417218 186348 417454
rect 186000 417134 186348 417218
rect 186000 416898 186056 417134
rect 186292 416898 186348 417134
rect 186000 416866 186348 416898
rect 45234 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 45854 406894
rect 45234 406574 45854 406658
rect 45234 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 45854 406574
rect 45234 370894 45854 406338
rect 50952 399454 51300 399486
rect 50952 399218 51008 399454
rect 51244 399218 51300 399454
rect 50952 399134 51300 399218
rect 50952 398898 51008 399134
rect 51244 398898 51300 399134
rect 50952 398866 51300 398898
rect 185320 399454 185668 399486
rect 185320 399218 185376 399454
rect 185612 399218 185668 399454
rect 185320 399134 185668 399218
rect 185320 398898 185376 399134
rect 185612 398898 185668 399134
rect 185320 398866 185668 398898
rect 50272 381454 50620 381486
rect 50272 381218 50328 381454
rect 50564 381218 50620 381454
rect 50272 381134 50620 381218
rect 50272 380898 50328 381134
rect 50564 380898 50620 381134
rect 50272 380866 50620 380898
rect 186000 381454 186348 381486
rect 186000 381218 186056 381454
rect 186292 381218 186348 381454
rect 186000 381134 186348 381218
rect 186000 380898 186056 381134
rect 186292 380898 186348 381134
rect 186000 380866 186348 380898
rect 66056 379810 66116 380106
rect 67144 379810 67204 380106
rect 68232 379810 68292 380106
rect 69592 379810 69652 380106
rect 70544 379810 70604 380106
rect 66056 379750 66178 379810
rect 67144 379750 67282 379810
rect 68232 379750 68386 379810
rect 69592 379750 69674 379810
rect 45234 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 45854 370894
rect 45234 370574 45854 370658
rect 45234 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 45854 370574
rect 45234 334894 45854 370338
rect 45234 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 45854 334894
rect 45234 334574 45854 334658
rect 45234 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 45854 334574
rect 45234 298894 45854 334338
rect 45234 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 45854 298894
rect 45234 298574 45854 298658
rect 45234 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 45854 298574
rect 45234 262894 45854 298338
rect 48954 374614 49574 378000
rect 48954 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 49574 374614
rect 48954 374294 49574 374378
rect 48954 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 49574 374294
rect 48954 338614 49574 374058
rect 48954 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 49574 338614
rect 48954 338294 49574 338378
rect 48954 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 49574 338294
rect 48954 302614 49574 338058
rect 48954 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 49574 302614
rect 48954 302294 49574 302378
rect 48954 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 49574 302294
rect 48954 285308 49574 302058
rect 55794 345454 56414 378000
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 285308 56414 308898
rect 59514 349174 60134 378000
rect 59514 348938 59546 349174
rect 59782 348938 59866 349174
rect 60102 348938 60134 349174
rect 59514 348854 60134 348938
rect 59514 348618 59546 348854
rect 59782 348618 59866 348854
rect 60102 348618 60134 348854
rect 59514 313174 60134 348618
rect 59514 312938 59546 313174
rect 59782 312938 59866 313174
rect 60102 312938 60134 313174
rect 59514 312854 60134 312938
rect 59514 312618 59546 312854
rect 59782 312618 59866 312854
rect 60102 312618 60134 312854
rect 59514 285308 60134 312618
rect 63234 352894 63854 378000
rect 66118 377093 66178 379750
rect 67222 378181 67282 379750
rect 67219 378180 67285 378181
rect 67219 378116 67220 378180
rect 67284 378116 67285 378180
rect 67219 378115 67285 378116
rect 66115 377092 66181 377093
rect 66115 377028 66116 377092
rect 66180 377028 66181 377092
rect 66115 377027 66181 377028
rect 63234 352658 63266 352894
rect 63502 352658 63586 352894
rect 63822 352658 63854 352894
rect 63234 352574 63854 352658
rect 63234 352338 63266 352574
rect 63502 352338 63586 352574
rect 63822 352338 63854 352574
rect 63234 316894 63854 352338
rect 63234 316658 63266 316894
rect 63502 316658 63586 316894
rect 63822 316658 63854 316894
rect 63234 316574 63854 316658
rect 63234 316338 63266 316574
rect 63502 316338 63586 316574
rect 63822 316338 63854 316574
rect 63234 285308 63854 316338
rect 66954 356614 67574 378000
rect 68326 377093 68386 379750
rect 69614 377093 69674 379750
rect 70534 379750 70604 379810
rect 71768 379810 71828 380106
rect 73128 379810 73188 380106
rect 74216 379810 74276 380106
rect 71768 379750 71882 379810
rect 70534 377093 70594 379750
rect 71822 377093 71882 379750
rect 73110 379750 73188 379810
rect 74214 379750 74276 379810
rect 75440 379810 75500 380106
rect 76528 379810 76588 380106
rect 77616 379810 77676 380106
rect 78296 379810 78356 380106
rect 75440 379750 75562 379810
rect 76528 379750 76666 379810
rect 77616 379750 77770 379810
rect 68323 377092 68389 377093
rect 68323 377028 68324 377092
rect 68388 377028 68389 377092
rect 68323 377027 68389 377028
rect 69611 377092 69677 377093
rect 69611 377028 69612 377092
rect 69676 377028 69677 377092
rect 69611 377027 69677 377028
rect 70531 377092 70597 377093
rect 70531 377028 70532 377092
rect 70596 377028 70597 377092
rect 70531 377027 70597 377028
rect 71819 377092 71885 377093
rect 71819 377028 71820 377092
rect 71884 377028 71885 377092
rect 71819 377027 71885 377028
rect 73110 376957 73170 379750
rect 74214 378181 74274 379750
rect 74211 378180 74277 378181
rect 74211 378116 74212 378180
rect 74276 378116 74277 378180
rect 74211 378115 74277 378116
rect 73107 376956 73173 376957
rect 73107 376892 73108 376956
rect 73172 376892 73173 376956
rect 73107 376891 73173 376892
rect 66954 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 67574 356614
rect 66954 356294 67574 356378
rect 66954 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 67574 356294
rect 66954 320614 67574 356058
rect 66954 320378 66986 320614
rect 67222 320378 67306 320614
rect 67542 320378 67574 320614
rect 66954 320294 67574 320378
rect 66954 320058 66986 320294
rect 67222 320058 67306 320294
rect 67542 320058 67574 320294
rect 66954 285308 67574 320058
rect 73794 363454 74414 378000
rect 75502 377093 75562 379750
rect 76606 377093 76666 379750
rect 77710 378181 77770 379750
rect 78262 379750 78356 379810
rect 78704 379810 78764 380106
rect 80064 379810 80124 380106
rect 80744 379810 80804 380106
rect 81288 379810 81348 380106
rect 78704 379750 78874 379810
rect 80064 379750 80162 379810
rect 80744 379750 80898 379810
rect 77707 378180 77773 378181
rect 77707 378116 77708 378180
rect 77772 378116 77773 378180
rect 77707 378115 77773 378116
rect 75499 377092 75565 377093
rect 75499 377028 75500 377092
rect 75564 377028 75565 377092
rect 75499 377027 75565 377028
rect 76603 377092 76669 377093
rect 76603 377028 76604 377092
rect 76668 377028 76669 377092
rect 76603 377027 76669 377028
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 73794 327454 74414 362898
rect 73794 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 74414 327454
rect 73794 327134 74414 327218
rect 73794 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 74414 327134
rect 73794 291454 74414 326898
rect 73794 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 74414 291454
rect 73794 291134 74414 291218
rect 73794 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 74414 291134
rect 73794 285308 74414 290898
rect 77514 367174 78134 378000
rect 78262 377093 78322 379750
rect 78814 377093 78874 379750
rect 80102 377093 80162 379750
rect 78259 377092 78325 377093
rect 78259 377028 78260 377092
rect 78324 377028 78325 377092
rect 78259 377027 78325 377028
rect 78811 377092 78877 377093
rect 78811 377028 78812 377092
rect 78876 377028 78877 377092
rect 78811 377027 78877 377028
rect 80099 377092 80165 377093
rect 80099 377028 80100 377092
rect 80164 377028 80165 377092
rect 80099 377027 80165 377028
rect 80838 376957 80898 379750
rect 81206 379750 81348 379810
rect 82376 379810 82436 380106
rect 83464 379810 83524 380106
rect 83600 379810 83660 380106
rect 82376 379750 82554 379810
rect 81206 378181 81266 379750
rect 81203 378180 81269 378181
rect 81203 378116 81204 378180
rect 81268 378116 81269 378180
rect 81203 378115 81269 378116
rect 80835 376956 80901 376957
rect 80835 376892 80836 376956
rect 80900 376892 80901 376956
rect 80835 376891 80901 376892
rect 77514 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 78134 367174
rect 77514 366854 78134 366938
rect 77514 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 78134 366854
rect 77514 331174 78134 366618
rect 77514 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 78134 331174
rect 77514 330854 78134 330938
rect 77514 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 78134 330854
rect 77514 295174 78134 330618
rect 77514 294938 77546 295174
rect 77782 294938 77866 295174
rect 78102 294938 78134 295174
rect 77514 294854 78134 294938
rect 77514 294618 77546 294854
rect 77782 294618 77866 294854
rect 78102 294618 78134 294854
rect 77514 285308 78134 294618
rect 81234 370894 81854 378000
rect 82494 377093 82554 379750
rect 83414 379750 83524 379810
rect 83598 379750 83660 379810
rect 82491 377092 82557 377093
rect 82491 377028 82492 377092
rect 82556 377028 82557 377092
rect 82491 377027 82557 377028
rect 83414 376957 83474 379750
rect 83598 377093 83658 379750
rect 84552 379530 84612 380106
rect 85912 379810 85972 380106
rect 84518 379470 84612 379530
rect 85806 379750 85972 379810
rect 84518 377093 84578 379470
rect 85806 378045 85866 379750
rect 86048 379530 86108 380106
rect 87000 379541 87060 380106
rect 88088 379541 88148 380106
rect 85990 379470 86108 379530
rect 86997 379540 87063 379541
rect 86997 379476 86998 379540
rect 87062 379476 87063 379540
rect 86997 379475 87063 379476
rect 88085 379540 88151 379541
rect 88085 379476 88086 379540
rect 88150 379476 88151 379540
rect 88085 379475 88151 379476
rect 88496 379530 88556 380106
rect 89448 379541 89508 380106
rect 90672 379541 90732 380106
rect 89445 379540 89511 379541
rect 88496 379470 88626 379530
rect 89445 379476 89446 379540
rect 89510 379476 89511 379540
rect 89445 379475 89511 379476
rect 90669 379540 90735 379541
rect 90669 379476 90670 379540
rect 90734 379476 90735 379540
rect 90669 379475 90735 379476
rect 91080 379530 91140 380106
rect 91760 379530 91820 380106
rect 92848 379530 92908 380106
rect 91080 379470 91202 379530
rect 91760 379470 91938 379530
rect 85803 378044 85869 378045
rect 83595 377092 83661 377093
rect 83595 377028 83596 377092
rect 83660 377028 83661 377092
rect 83595 377027 83661 377028
rect 84515 377092 84581 377093
rect 84515 377028 84516 377092
rect 84580 377028 84581 377092
rect 84515 377027 84581 377028
rect 83411 376956 83477 376957
rect 83411 376892 83412 376956
rect 83476 376892 83477 376956
rect 83411 376891 83477 376892
rect 81234 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 81854 370894
rect 81234 370574 81854 370658
rect 81234 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 81854 370574
rect 81234 334894 81854 370338
rect 81234 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 81854 334894
rect 81234 334574 81854 334658
rect 81234 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 81854 334574
rect 81234 298894 81854 334338
rect 81234 298658 81266 298894
rect 81502 298658 81586 298894
rect 81822 298658 81854 298894
rect 81234 298574 81854 298658
rect 81234 298338 81266 298574
rect 81502 298338 81586 298574
rect 81822 298338 81854 298574
rect 78811 285700 78877 285701
rect 78811 285636 78812 285700
rect 78876 285636 78877 285700
rect 78811 285635 78877 285636
rect 81019 285700 81085 285701
rect 81019 285636 81020 285700
rect 81084 285636 81085 285700
rect 81019 285635 81085 285636
rect 78814 283930 78874 285635
rect 81022 283930 81082 285635
rect 81234 285308 81854 298338
rect 84954 374614 85574 378000
rect 85803 377980 85804 378044
rect 85868 377980 85869 378044
rect 85803 377979 85869 377980
rect 85990 377093 86050 379470
rect 88566 377093 88626 379470
rect 91142 377093 91202 379470
rect 91878 378181 91938 379470
rect 92798 379470 92908 379530
rect 93528 379530 93588 380106
rect 93936 379530 93996 380106
rect 95296 379530 95356 380106
rect 95976 379530 96036 380106
rect 93528 379470 93594 379530
rect 91875 378180 91941 378181
rect 91875 378116 91876 378180
rect 91940 378116 91941 378180
rect 91875 378115 91941 378116
rect 92798 378045 92858 379470
rect 92795 378044 92861 378045
rect 85987 377092 86053 377093
rect 85987 377028 85988 377092
rect 86052 377028 86053 377092
rect 85987 377027 86053 377028
rect 88563 377092 88629 377093
rect 88563 377028 88564 377092
rect 88628 377028 88629 377092
rect 88563 377027 88629 377028
rect 91139 377092 91205 377093
rect 91139 377028 91140 377092
rect 91204 377028 91205 377092
rect 91139 377027 91205 377028
rect 84954 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 85574 374614
rect 84954 374294 85574 374378
rect 84954 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 85574 374294
rect 84954 338614 85574 374058
rect 84954 338378 84986 338614
rect 85222 338378 85306 338614
rect 85542 338378 85574 338614
rect 84954 338294 85574 338378
rect 84954 338058 84986 338294
rect 85222 338058 85306 338294
rect 85542 338058 85574 338294
rect 84954 302614 85574 338058
rect 84954 302378 84986 302614
rect 85222 302378 85306 302614
rect 85542 302378 85574 302614
rect 84954 302294 85574 302378
rect 84954 302058 84986 302294
rect 85222 302058 85306 302294
rect 85542 302058 85574 302294
rect 83411 285700 83477 285701
rect 83411 285636 83412 285700
rect 83476 285636 83477 285700
rect 83411 285635 83477 285636
rect 78704 283870 78874 283930
rect 81016 283870 81082 283930
rect 83414 283930 83474 285635
rect 84954 285308 85574 302058
rect 91794 345454 92414 378000
rect 92795 377980 92796 378044
rect 92860 377980 92861 378044
rect 92795 377979 92861 377980
rect 93534 377093 93594 379470
rect 93902 379470 93996 379530
rect 95190 379470 95356 379530
rect 95926 379470 96036 379530
rect 96384 379530 96444 380106
rect 97608 379530 97668 380106
rect 96384 379470 96538 379530
rect 93902 378045 93962 379470
rect 95190 378045 95250 379470
rect 95926 378181 95986 379470
rect 95923 378180 95989 378181
rect 95923 378116 95924 378180
rect 95988 378116 95989 378180
rect 95923 378115 95989 378116
rect 93899 378044 93965 378045
rect 93899 377980 93900 378044
rect 93964 377980 93965 378044
rect 93899 377979 93965 377980
rect 95187 378044 95253 378045
rect 95187 377980 95188 378044
rect 95252 377980 95253 378044
rect 95187 377979 95253 377980
rect 93531 377092 93597 377093
rect 93531 377028 93532 377092
rect 93596 377028 93597 377092
rect 93531 377027 93597 377028
rect 91794 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 92414 345454
rect 91794 345134 92414 345218
rect 91794 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 92414 345134
rect 91794 309454 92414 344898
rect 91794 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 92414 309454
rect 91794 309134 92414 309218
rect 91794 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 92414 309134
rect 86171 285700 86237 285701
rect 86171 285636 86172 285700
rect 86236 285636 86237 285700
rect 86171 285635 86237 285636
rect 88563 285700 88629 285701
rect 88563 285636 88564 285700
rect 88628 285636 88629 285700
rect 88563 285635 88629 285636
rect 86174 283930 86234 285635
rect 88566 283930 88626 285635
rect 91794 285308 92414 308898
rect 95514 349174 96134 378000
rect 96478 377909 96538 379470
rect 97582 379470 97668 379530
rect 98288 379530 98348 380106
rect 98696 379530 98756 380106
rect 98288 379470 98378 379530
rect 97582 378045 97642 379470
rect 97579 378044 97645 378045
rect 97579 377980 97580 378044
rect 97644 377980 97645 378044
rect 97579 377979 97645 377980
rect 96475 377908 96541 377909
rect 96475 377844 96476 377908
rect 96540 377844 96541 377908
rect 96475 377843 96541 377844
rect 98318 377093 98378 379470
rect 98686 379470 98756 379530
rect 99784 379530 99844 380106
rect 101008 379530 101068 380106
rect 101144 379810 101204 380106
rect 101144 379750 101322 379810
rect 99784 379470 99850 379530
rect 101008 379470 101138 379530
rect 98686 378997 98746 379470
rect 98683 378996 98749 378997
rect 98683 378932 98684 378996
rect 98748 378932 98749 378996
rect 98683 378931 98749 378932
rect 99790 378181 99850 379470
rect 99787 378180 99853 378181
rect 99787 378116 99788 378180
rect 99852 378116 99853 378180
rect 99787 378115 99853 378116
rect 98315 377092 98381 377093
rect 98315 377028 98316 377092
rect 98380 377028 98381 377092
rect 98315 377027 98381 377028
rect 95514 348938 95546 349174
rect 95782 348938 95866 349174
rect 96102 348938 96134 349174
rect 95514 348854 96134 348938
rect 95514 348618 95546 348854
rect 95782 348618 95866 348854
rect 96102 348618 96134 348854
rect 95514 313174 96134 348618
rect 95514 312938 95546 313174
rect 95782 312938 95866 313174
rect 96102 312938 96134 313174
rect 95514 312854 96134 312938
rect 95514 312618 95546 312854
rect 95782 312618 95866 312854
rect 96102 312618 96134 312854
rect 93531 285700 93597 285701
rect 93531 285636 93532 285700
rect 93596 285636 93597 285700
rect 93531 285635 93597 285636
rect 91139 284884 91205 284885
rect 91139 284820 91140 284884
rect 91204 284820 91205 284884
rect 91139 284819 91205 284820
rect 91142 283930 91202 284819
rect 93534 283930 93594 285635
rect 95514 285308 96134 312618
rect 99234 352894 99854 378000
rect 101078 377773 101138 379470
rect 101262 379405 101322 379750
rect 102232 379530 102292 380106
rect 103320 379810 103380 380106
rect 102182 379470 102292 379530
rect 103286 379750 103380 379810
rect 101259 379404 101325 379405
rect 101259 379340 101260 379404
rect 101324 379340 101325 379404
rect 101259 379339 101325 379340
rect 101075 377772 101141 377773
rect 101075 377708 101076 377772
rect 101140 377708 101141 377772
rect 101075 377707 101141 377708
rect 102182 377093 102242 379470
rect 103286 379269 103346 379750
rect 103592 379674 103652 380106
rect 104408 379674 104468 380106
rect 105768 379810 105828 380106
rect 105768 379750 105922 379810
rect 103592 379614 103714 379674
rect 103283 379268 103349 379269
rect 103283 379204 103284 379268
rect 103348 379204 103349 379268
rect 103283 379203 103349 379204
rect 103654 378181 103714 379614
rect 104390 379614 104468 379674
rect 103651 378180 103717 378181
rect 103651 378116 103652 378180
rect 103716 378116 103717 378180
rect 103651 378115 103717 378116
rect 102179 377092 102245 377093
rect 102179 377028 102180 377092
rect 102244 377028 102245 377092
rect 102179 377027 102245 377028
rect 99234 352658 99266 352894
rect 99502 352658 99586 352894
rect 99822 352658 99854 352894
rect 99234 352574 99854 352658
rect 99234 352338 99266 352574
rect 99502 352338 99586 352574
rect 99822 352338 99854 352574
rect 99234 316894 99854 352338
rect 99234 316658 99266 316894
rect 99502 316658 99586 316894
rect 99822 316658 99854 316894
rect 99234 316574 99854 316658
rect 99234 316338 99266 316574
rect 99502 316338 99586 316574
rect 99822 316338 99854 316574
rect 99234 285308 99854 316338
rect 102954 356614 103574 378000
rect 104390 377909 104450 379614
rect 104387 377908 104453 377909
rect 104387 377844 104388 377908
rect 104452 377844 104453 377908
rect 104387 377843 104453 377844
rect 105862 377501 105922 379750
rect 106040 379674 106100 380106
rect 106992 379674 107052 380106
rect 108080 379674 108140 380106
rect 108488 379674 108548 380106
rect 106040 379614 106106 379674
rect 106046 378045 106106 379614
rect 106966 379614 107052 379674
rect 108070 379614 108140 379674
rect 108438 379614 108548 379674
rect 109168 379674 109228 380106
rect 110936 379677 110996 380106
rect 113520 379677 113580 380106
rect 115968 379810 116028 380106
rect 115968 379750 116042 379810
rect 110933 379676 110999 379677
rect 109168 379614 109234 379674
rect 106043 378044 106109 378045
rect 106043 377980 106044 378044
rect 106108 377980 106109 378044
rect 106043 377979 106109 377980
rect 106966 377773 107026 379614
rect 106963 377772 107029 377773
rect 106963 377708 106964 377772
rect 107028 377708 107029 377772
rect 106963 377707 107029 377708
rect 108070 377637 108130 379614
rect 108438 378045 108498 379614
rect 109174 379133 109234 379614
rect 110933 379612 110934 379676
rect 110998 379612 110999 379676
rect 110933 379611 110999 379612
rect 113517 379676 113583 379677
rect 113517 379612 113518 379676
rect 113582 379612 113583 379676
rect 113517 379611 113583 379612
rect 115982 379541 116042 379750
rect 118280 379677 118340 380106
rect 121000 379677 121060 380106
rect 123448 379677 123508 380106
rect 125896 379810 125956 380106
rect 128480 379810 128540 380106
rect 125896 379750 125978 379810
rect 128480 379750 128554 379810
rect 118277 379676 118343 379677
rect 118277 379612 118278 379676
rect 118342 379612 118343 379676
rect 118277 379611 118343 379612
rect 120997 379676 121063 379677
rect 120997 379612 120998 379676
rect 121062 379612 121063 379676
rect 120997 379611 121063 379612
rect 123445 379676 123511 379677
rect 123445 379612 123446 379676
rect 123510 379612 123511 379676
rect 123445 379611 123511 379612
rect 115979 379540 116045 379541
rect 115979 379476 115980 379540
rect 116044 379476 116045 379540
rect 115979 379475 116045 379476
rect 109171 379132 109237 379133
rect 109171 379068 109172 379132
rect 109236 379068 109237 379132
rect 109171 379067 109237 379068
rect 125918 378045 125978 379750
rect 128494 378181 128554 379750
rect 130928 379677 130988 380106
rect 133512 379810 133572 380106
rect 133462 379750 133572 379810
rect 135960 379810 136020 380106
rect 138544 379810 138604 380106
rect 140992 379810 141052 380106
rect 135960 379750 136098 379810
rect 138544 379750 138674 379810
rect 140992 379750 141066 379810
rect 130925 379676 130991 379677
rect 130925 379612 130926 379676
rect 130990 379612 130991 379676
rect 130925 379611 130991 379612
rect 128491 378180 128557 378181
rect 128491 378116 128492 378180
rect 128556 378116 128557 378180
rect 128491 378115 128557 378116
rect 133462 378045 133522 379750
rect 136038 378045 136098 379750
rect 138614 378045 138674 379750
rect 141006 378045 141066 379750
rect 143440 379677 143500 380106
rect 145888 379810 145948 380106
rect 148472 379810 148532 380106
rect 150920 379810 150980 380106
rect 153368 379810 153428 380106
rect 155952 379810 156012 380106
rect 173224 379810 173284 380106
rect 145888 379750 146034 379810
rect 148472 379750 148610 379810
rect 150920 379750 151002 379810
rect 143437 379676 143503 379677
rect 143437 379612 143438 379676
rect 143502 379612 143503 379676
rect 143437 379611 143503 379612
rect 145974 378181 146034 379750
rect 145971 378180 146037 378181
rect 145971 378116 145972 378180
rect 146036 378116 146037 378180
rect 145971 378115 146037 378116
rect 148550 378045 148610 379750
rect 150942 379541 151002 379750
rect 153334 379750 153428 379810
rect 155910 379750 156012 379810
rect 173206 379750 173284 379810
rect 173360 379810 173420 380106
rect 173360 379750 173450 379810
rect 150939 379540 151005 379541
rect 150939 379476 150940 379540
rect 151004 379476 151005 379540
rect 150939 379475 151005 379476
rect 153334 378181 153394 379750
rect 153331 378180 153397 378181
rect 153331 378116 153332 378180
rect 153396 378116 153397 378180
rect 153331 378115 153397 378116
rect 155910 378045 155970 379750
rect 108435 378044 108501 378045
rect 108435 377980 108436 378044
rect 108500 377980 108501 378044
rect 125915 378044 125981 378045
rect 108435 377979 108501 377980
rect 108067 377636 108133 377637
rect 108067 377572 108068 377636
rect 108132 377572 108133 377636
rect 108067 377571 108133 377572
rect 105859 377500 105925 377501
rect 105859 377436 105860 377500
rect 105924 377436 105925 377500
rect 105859 377435 105925 377436
rect 102954 356378 102986 356614
rect 103222 356378 103306 356614
rect 103542 356378 103574 356614
rect 102954 356294 103574 356378
rect 102954 356058 102986 356294
rect 103222 356058 103306 356294
rect 103542 356058 103574 356294
rect 102954 320614 103574 356058
rect 102954 320378 102986 320614
rect 103222 320378 103306 320614
rect 103542 320378 103574 320614
rect 102954 320294 103574 320378
rect 102954 320058 102986 320294
rect 103222 320058 103306 320294
rect 103542 320058 103574 320294
rect 101259 285700 101325 285701
rect 101259 285636 101260 285700
rect 101324 285636 101325 285700
rect 101259 285635 101325 285636
rect 96107 285156 96173 285157
rect 96107 285092 96108 285156
rect 96172 285092 96173 285156
rect 96107 285091 96173 285092
rect 83414 283870 83524 283930
rect 86174 283870 86244 283930
rect 78704 283220 78764 283870
rect 81016 283220 81076 283870
rect 83464 283220 83524 283870
rect 86184 283220 86244 283870
rect 88496 283870 88626 283930
rect 91080 283870 91202 283930
rect 93528 283870 93594 283930
rect 96110 283930 96170 285091
rect 98499 285020 98565 285021
rect 98499 284956 98500 285020
rect 98564 284956 98565 285020
rect 98499 284955 98565 284956
rect 98502 283930 98562 284955
rect 101262 283930 101322 285635
rect 102954 285308 103574 320058
rect 109794 363454 110414 378000
rect 109794 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 110414 363454
rect 109794 363134 110414 363218
rect 109794 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 110414 363134
rect 109794 327454 110414 362898
rect 109794 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 110414 327454
rect 109794 327134 110414 327218
rect 109794 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 110414 327134
rect 109794 291454 110414 326898
rect 109794 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 110414 291454
rect 109794 291134 110414 291218
rect 109794 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 110414 291134
rect 108435 285972 108501 285973
rect 108435 285908 108436 285972
rect 108500 285908 108501 285972
rect 108435 285907 108501 285908
rect 103835 285700 103901 285701
rect 103835 285636 103836 285700
rect 103900 285636 103901 285700
rect 103835 285635 103901 285636
rect 106227 285700 106293 285701
rect 106227 285636 106228 285700
rect 106292 285636 106293 285700
rect 106227 285635 106293 285636
rect 103838 283930 103898 285635
rect 106230 283930 106290 285635
rect 96110 283870 96172 283930
rect 98502 283870 98620 283930
rect 88496 283220 88556 283870
rect 91080 283220 91140 283870
rect 93528 283220 93588 283870
rect 96112 283220 96172 283870
rect 98560 283220 98620 283870
rect 101144 283870 101322 283930
rect 103592 283870 103898 283930
rect 106176 283870 106290 283930
rect 108438 283930 108498 285907
rect 109794 285308 110414 290898
rect 113514 367174 114134 378000
rect 113514 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 114134 367174
rect 113514 366854 114134 366938
rect 113514 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 114134 366854
rect 113514 331174 114134 366618
rect 113514 330938 113546 331174
rect 113782 330938 113866 331174
rect 114102 330938 114134 331174
rect 113514 330854 114134 330938
rect 113514 330618 113546 330854
rect 113782 330618 113866 330854
rect 114102 330618 114134 330854
rect 113514 295174 114134 330618
rect 113514 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 114134 295174
rect 113514 294854 114134 294938
rect 113514 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 114134 294854
rect 111011 285972 111077 285973
rect 111011 285908 111012 285972
rect 111076 285908 111077 285972
rect 111011 285907 111077 285908
rect 111014 283930 111074 285907
rect 113514 285308 114134 294618
rect 117234 370894 117854 378000
rect 117234 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 117854 370894
rect 117234 370574 117854 370658
rect 117234 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 117854 370574
rect 117234 334894 117854 370338
rect 117234 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 117854 334894
rect 117234 334574 117854 334658
rect 117234 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 117854 334574
rect 117234 298894 117854 334338
rect 117234 298658 117266 298894
rect 117502 298658 117586 298894
rect 117822 298658 117854 298894
rect 117234 298574 117854 298658
rect 117234 298338 117266 298574
rect 117502 298338 117586 298574
rect 117822 298338 117854 298574
rect 116163 286516 116229 286517
rect 116163 286452 116164 286516
rect 116228 286452 116229 286516
rect 116163 286451 116229 286452
rect 113771 285156 113837 285157
rect 113771 285092 113772 285156
rect 113836 285092 113837 285156
rect 113771 285091 113837 285092
rect 113774 283930 113834 285091
rect 116166 283930 116226 286451
rect 117234 285308 117854 298338
rect 120954 374614 121574 378000
rect 125915 377980 125916 378044
rect 125980 377980 125981 378044
rect 133459 378044 133525 378045
rect 125915 377979 125981 377980
rect 120954 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 121574 374614
rect 120954 374294 121574 374378
rect 120954 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 121574 374294
rect 120954 338614 121574 374058
rect 120954 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 121574 338614
rect 120954 338294 121574 338378
rect 120954 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 121574 338294
rect 120954 302614 121574 338058
rect 120954 302378 120986 302614
rect 121222 302378 121306 302614
rect 121542 302378 121574 302614
rect 120954 302294 121574 302378
rect 120954 302058 120986 302294
rect 121222 302058 121306 302294
rect 121542 302058 121574 302294
rect 120763 285700 120829 285701
rect 120763 285636 120764 285700
rect 120828 285636 120829 285700
rect 120763 285635 120829 285636
rect 118555 285020 118621 285021
rect 118555 284956 118556 285020
rect 118620 284956 118621 285020
rect 118555 284955 118621 284956
rect 118558 283930 118618 284955
rect 108438 283870 108548 283930
rect 101144 283220 101204 283870
rect 103592 283220 103652 283870
rect 106176 283220 106236 283870
rect 108488 283220 108548 283870
rect 110936 283870 111074 283930
rect 113656 283870 113834 283930
rect 116104 283870 116226 283930
rect 118552 283870 118618 283930
rect 120766 283930 120826 285635
rect 120954 285308 121574 302058
rect 127794 345454 128414 378000
rect 127794 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 128414 345454
rect 127794 345134 128414 345218
rect 127794 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 128414 345134
rect 127794 309454 128414 344898
rect 127794 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 128414 309454
rect 127794 309134 128414 309218
rect 127794 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 128414 309134
rect 125915 286108 125981 286109
rect 125915 286044 125916 286108
rect 125980 286044 125981 286108
rect 125915 286043 125981 286044
rect 123523 285156 123589 285157
rect 123523 285092 123524 285156
rect 123588 285092 123589 285156
rect 123523 285091 123589 285092
rect 123526 283930 123586 285091
rect 125918 283930 125978 286043
rect 127794 285308 128414 308898
rect 131514 349174 132134 378000
rect 133459 377980 133460 378044
rect 133524 377980 133525 378044
rect 136035 378044 136101 378045
rect 133459 377979 133525 377980
rect 131514 348938 131546 349174
rect 131782 348938 131866 349174
rect 132102 348938 132134 349174
rect 131514 348854 132134 348938
rect 131514 348618 131546 348854
rect 131782 348618 131866 348854
rect 132102 348618 132134 348854
rect 131514 313174 132134 348618
rect 131514 312938 131546 313174
rect 131782 312938 131866 313174
rect 132102 312938 132134 313174
rect 131514 312854 132134 312938
rect 131514 312618 131546 312854
rect 131782 312618 131866 312854
rect 132102 312618 132134 312854
rect 131067 286108 131133 286109
rect 131067 286044 131068 286108
rect 131132 286044 131133 286108
rect 131067 286043 131133 286044
rect 128675 285156 128741 285157
rect 128675 285092 128676 285156
rect 128740 285092 128741 285156
rect 128675 285091 128741 285092
rect 128678 283930 128738 285091
rect 131070 283930 131130 286043
rect 131514 285308 132134 312618
rect 135234 352894 135854 378000
rect 136035 377980 136036 378044
rect 136100 377980 136101 378044
rect 136035 377979 136101 377980
rect 138611 378044 138677 378045
rect 138611 377980 138612 378044
rect 138676 377980 138677 378044
rect 141003 378044 141069 378045
rect 138611 377979 138677 377980
rect 135234 352658 135266 352894
rect 135502 352658 135586 352894
rect 135822 352658 135854 352894
rect 135234 352574 135854 352658
rect 135234 352338 135266 352574
rect 135502 352338 135586 352574
rect 135822 352338 135854 352574
rect 135234 316894 135854 352338
rect 135234 316658 135266 316894
rect 135502 316658 135586 316894
rect 135822 316658 135854 316894
rect 135234 316574 135854 316658
rect 135234 316338 135266 316574
rect 135502 316338 135586 316574
rect 135822 316338 135854 316574
rect 133459 286108 133525 286109
rect 133459 286044 133460 286108
rect 133524 286044 133525 286108
rect 133459 286043 133525 286044
rect 120766 283870 121060 283930
rect 123526 283870 123644 283930
rect 110936 283220 110996 283870
rect 113656 283220 113716 283870
rect 116104 283220 116164 283870
rect 118552 283220 118612 283870
rect 121000 283220 121060 283870
rect 123584 283220 123644 283870
rect 125896 283870 125978 283930
rect 128616 283870 128738 283930
rect 131064 283870 131130 283930
rect 133462 283930 133522 286043
rect 135234 285308 135854 316338
rect 138954 356614 139574 378000
rect 141003 377980 141004 378044
rect 141068 377980 141069 378044
rect 148547 378044 148613 378045
rect 141003 377979 141069 377980
rect 138954 356378 138986 356614
rect 139222 356378 139306 356614
rect 139542 356378 139574 356614
rect 138954 356294 139574 356378
rect 138954 356058 138986 356294
rect 139222 356058 139306 356294
rect 139542 356058 139574 356294
rect 138954 320614 139574 356058
rect 138954 320378 138986 320614
rect 139222 320378 139306 320614
rect 139542 320378 139574 320614
rect 138954 320294 139574 320378
rect 138954 320058 138986 320294
rect 139222 320058 139306 320294
rect 139542 320058 139574 320294
rect 136035 286380 136101 286381
rect 136035 286316 136036 286380
rect 136100 286316 136101 286380
rect 136035 286315 136101 286316
rect 136038 283930 136098 286315
rect 138427 285700 138493 285701
rect 138427 285636 138428 285700
rect 138492 285636 138493 285700
rect 138427 285635 138493 285636
rect 138430 283930 138490 285635
rect 138954 285308 139574 320058
rect 145794 363454 146414 378000
rect 148547 377980 148548 378044
rect 148612 377980 148613 378044
rect 155907 378044 155973 378045
rect 148547 377979 148613 377980
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 145794 327454 146414 362898
rect 145794 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 146414 327454
rect 145794 327134 146414 327218
rect 145794 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 146414 327134
rect 145794 291454 146414 326898
rect 145794 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 146414 291454
rect 145794 291134 146414 291218
rect 145794 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 146414 291134
rect 141003 285700 141069 285701
rect 141003 285636 141004 285700
rect 141068 285636 141069 285700
rect 141003 285635 141069 285636
rect 143579 285700 143645 285701
rect 143579 285636 143580 285700
rect 143644 285636 143645 285700
rect 143579 285635 143645 285636
rect 145603 285700 145669 285701
rect 145603 285636 145604 285700
rect 145668 285636 145669 285700
rect 145603 285635 145669 285636
rect 141006 283930 141066 285635
rect 143582 283930 143642 285635
rect 133462 283870 133572 283930
rect 125896 283220 125956 283870
rect 128616 283220 128676 283870
rect 131064 283220 131124 283870
rect 133512 283220 133572 283870
rect 135960 283870 136098 283930
rect 138408 283870 138490 283930
rect 140992 283870 141066 283930
rect 143576 283870 143642 283930
rect 145606 283930 145666 285635
rect 145794 285308 146414 290898
rect 149514 367174 150134 378000
rect 149514 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 150134 367174
rect 149514 366854 150134 366938
rect 149514 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 150134 366854
rect 149514 331174 150134 366618
rect 149514 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 150134 331174
rect 149514 330854 150134 330938
rect 149514 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 150134 330854
rect 149514 295174 150134 330618
rect 149514 294938 149546 295174
rect 149782 294938 149866 295174
rect 150102 294938 150134 295174
rect 149514 294854 150134 294938
rect 149514 294618 149546 294854
rect 149782 294618 149866 294854
rect 150102 294618 150134 294854
rect 148547 285700 148613 285701
rect 148547 285636 148548 285700
rect 148612 285636 148613 285700
rect 148547 285635 148613 285636
rect 148550 283930 148610 285635
rect 149514 285308 150134 294618
rect 153234 370894 153854 378000
rect 155907 377980 155908 378044
rect 155972 377980 155973 378044
rect 155907 377979 155973 377980
rect 153234 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 153854 370894
rect 153234 370574 153854 370658
rect 153234 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 153854 370574
rect 153234 334894 153854 370338
rect 153234 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 153854 334894
rect 153234 334574 153854 334658
rect 153234 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 153854 334574
rect 153234 298894 153854 334338
rect 153234 298658 153266 298894
rect 153502 298658 153586 298894
rect 153822 298658 153854 298894
rect 153234 298574 153854 298658
rect 153234 298338 153266 298574
rect 153502 298338 153586 298574
rect 153822 298338 153854 298574
rect 151123 285700 151189 285701
rect 151123 285636 151124 285700
rect 151188 285636 151189 285700
rect 151123 285635 151189 285636
rect 151126 283930 151186 285635
rect 153234 285308 153854 298338
rect 156954 374614 157574 378000
rect 156954 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 157574 374614
rect 156954 374294 157574 374378
rect 156954 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 157574 374294
rect 156954 338614 157574 374058
rect 156954 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 157574 338614
rect 156954 338294 157574 338378
rect 156954 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 157574 338294
rect 156954 302614 157574 338058
rect 156954 302378 156986 302614
rect 157222 302378 157306 302614
rect 157542 302378 157574 302614
rect 156954 302294 157574 302378
rect 156954 302058 156986 302294
rect 157222 302058 157306 302294
rect 157542 302058 157574 302294
rect 154067 285700 154133 285701
rect 154067 285636 154068 285700
rect 154132 285636 154133 285700
rect 154067 285635 154133 285636
rect 156091 285700 156157 285701
rect 156091 285636 156092 285700
rect 156156 285636 156157 285700
rect 156091 285635 156157 285636
rect 154070 283930 154130 285635
rect 156094 283930 156154 285635
rect 156954 285308 157574 302058
rect 163794 345454 164414 378000
rect 163794 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 164414 345454
rect 163794 345134 164414 345218
rect 163794 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 164414 345134
rect 163794 309454 164414 344898
rect 163794 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 164414 309454
rect 163794 309134 164414 309218
rect 163794 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 164414 309134
rect 163794 285308 164414 308898
rect 167514 349174 168134 378000
rect 167514 348938 167546 349174
rect 167782 348938 167866 349174
rect 168102 348938 168134 349174
rect 167514 348854 168134 348938
rect 167514 348618 167546 348854
rect 167782 348618 167866 348854
rect 168102 348618 168134 348854
rect 167514 313174 168134 348618
rect 167514 312938 167546 313174
rect 167782 312938 167866 313174
rect 168102 312938 168134 313174
rect 167514 312854 168134 312938
rect 167514 312618 167546 312854
rect 167782 312618 167866 312854
rect 168102 312618 168134 312854
rect 167514 285308 168134 312618
rect 171234 352894 171854 378000
rect 173206 377229 173266 379750
rect 173203 377228 173269 377229
rect 173203 377164 173204 377228
rect 173268 377164 173269 377228
rect 173203 377163 173269 377164
rect 173390 376957 173450 379750
rect 173387 376956 173453 376957
rect 173387 376892 173388 376956
rect 173452 376892 173453 376956
rect 173387 376891 173453 376892
rect 171234 352658 171266 352894
rect 171502 352658 171586 352894
rect 171822 352658 171854 352894
rect 171234 352574 171854 352658
rect 171234 352338 171266 352574
rect 171502 352338 171586 352574
rect 171822 352338 171854 352574
rect 171234 316894 171854 352338
rect 171234 316658 171266 316894
rect 171502 316658 171586 316894
rect 171822 316658 171854 316894
rect 171234 316574 171854 316658
rect 171234 316338 171266 316574
rect 171502 316338 171586 316574
rect 171822 316338 171854 316574
rect 169707 286380 169773 286381
rect 169707 286316 169708 286380
rect 169772 286316 169773 286380
rect 169707 286315 169773 286316
rect 168419 286244 168485 286245
rect 168419 286180 168420 286244
rect 168484 286180 168485 286244
rect 168419 286179 168485 286180
rect 145606 283870 146084 283930
rect 135960 283220 136020 283870
rect 138408 283220 138468 283870
rect 140992 283220 141052 283870
rect 143576 283220 143636 283870
rect 146024 283220 146084 283870
rect 148472 283870 148610 283930
rect 151056 283870 151186 283930
rect 153368 283870 154130 283930
rect 156088 283870 156154 283930
rect 168422 283930 168482 286179
rect 169710 283930 169770 286315
rect 171234 285308 171854 316338
rect 174954 356614 175574 378000
rect 174954 356378 174986 356614
rect 175222 356378 175306 356614
rect 175542 356378 175574 356614
rect 174954 356294 175574 356378
rect 174954 356058 174986 356294
rect 175222 356058 175306 356294
rect 175542 356058 175574 356294
rect 174954 320614 175574 356058
rect 174954 320378 174986 320614
rect 175222 320378 175306 320614
rect 175542 320378 175574 320614
rect 174954 320294 175574 320378
rect 174954 320058 174986 320294
rect 175222 320058 175306 320294
rect 175542 320058 175574 320294
rect 174954 285308 175574 320058
rect 181794 363454 182414 378000
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 181794 327454 182414 362898
rect 181794 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 182414 327454
rect 181794 327134 182414 327218
rect 181794 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 182414 327134
rect 181794 291454 182414 326898
rect 181794 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 182414 291454
rect 181794 291134 182414 291218
rect 181794 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 182414 291134
rect 181794 285308 182414 290898
rect 185514 367174 186134 378000
rect 186822 377501 186882 460939
rect 186819 377500 186885 377501
rect 186819 377436 186820 377500
rect 186884 377436 186885 377500
rect 186819 377435 186885 377436
rect 187742 377365 187802 465155
rect 187739 377364 187805 377365
rect 187739 377300 187740 377364
rect 187804 377300 187805 377364
rect 187739 377299 187805 377300
rect 185514 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 186134 367174
rect 185514 366854 186134 366938
rect 185514 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 186134 366854
rect 185514 331174 186134 366618
rect 185514 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 186134 331174
rect 185514 330854 186134 330938
rect 185514 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 186134 330854
rect 185514 295174 186134 330618
rect 188294 317525 188354 465291
rect 189234 442894 189854 478338
rect 189234 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 189854 442894
rect 189234 442574 189854 442658
rect 189234 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 189854 442574
rect 189234 406894 189854 442338
rect 189234 406658 189266 406894
rect 189502 406658 189586 406894
rect 189822 406658 189854 406894
rect 189234 406574 189854 406658
rect 189234 406338 189266 406574
rect 189502 406338 189586 406574
rect 189822 406338 189854 406574
rect 189234 370894 189854 406338
rect 189234 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 189854 370894
rect 189234 370574 189854 370658
rect 189234 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 189854 370574
rect 189234 334894 189854 370338
rect 189234 334658 189266 334894
rect 189502 334658 189586 334894
rect 189822 334658 189854 334894
rect 189234 334574 189854 334658
rect 189234 334338 189266 334574
rect 189502 334338 189586 334574
rect 189822 334338 189854 334574
rect 188291 317524 188357 317525
rect 188291 317460 188292 317524
rect 188356 317460 188357 317524
rect 188291 317459 188357 317460
rect 185514 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 186134 295174
rect 185514 294854 186134 294938
rect 185514 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 186134 294854
rect 185514 285308 186134 294618
rect 189234 298894 189854 334338
rect 189234 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 189854 298894
rect 189234 298574 189854 298658
rect 189234 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 189854 298574
rect 188291 285836 188357 285837
rect 188291 285772 188292 285836
rect 188356 285772 188357 285836
rect 188291 285771 188357 285772
rect 180747 284068 180813 284069
rect 180747 284004 180748 284068
rect 180812 284004 180813 284068
rect 180747 284003 180813 284004
rect 168422 283870 168524 283930
rect 148472 283220 148532 283870
rect 151056 283220 151116 283870
rect 153368 283220 153428 283870
rect 156088 283220 156148 283870
rect 168464 283220 168524 283870
rect 169688 283870 169770 283930
rect 180750 283930 180810 284003
rect 180750 283870 180900 283930
rect 169688 283220 169748 283870
rect 180840 283220 180900 283870
rect 50272 273454 50620 273486
rect 50272 273218 50328 273454
rect 50564 273218 50620 273454
rect 50272 273134 50620 273218
rect 50272 272898 50328 273134
rect 50564 272898 50620 273134
rect 50272 272866 50620 272898
rect 186000 273454 186348 273486
rect 186000 273218 186056 273454
rect 186292 273218 186348 273454
rect 186000 273134 186348 273218
rect 186000 272898 186056 273134
rect 186292 272898 186348 273134
rect 186000 272866 186348 272898
rect 186819 270604 186885 270605
rect 186819 270540 186820 270604
rect 186884 270540 186885 270604
rect 186819 270539 186885 270540
rect 45234 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 45854 262894
rect 45234 262574 45854 262658
rect 45234 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 45854 262574
rect 45234 226894 45854 262338
rect 50952 255454 51300 255486
rect 50952 255218 51008 255454
rect 51244 255218 51300 255454
rect 50952 255134 51300 255218
rect 50952 254898 51008 255134
rect 51244 254898 51300 255134
rect 50952 254866 51300 254898
rect 185320 255454 185668 255486
rect 185320 255218 185376 255454
rect 185612 255218 185668 255454
rect 185320 255134 185668 255218
rect 185320 254898 185376 255134
rect 185612 254898 185668 255134
rect 185320 254866 185668 254898
rect 50272 237454 50620 237486
rect 50272 237218 50328 237454
rect 50564 237218 50620 237454
rect 50272 237134 50620 237218
rect 50272 236898 50328 237134
rect 50564 236898 50620 237134
rect 50272 236866 50620 236898
rect 186000 237454 186348 237486
rect 186000 237218 186056 237454
rect 186292 237218 186348 237454
rect 186000 237134 186348 237218
rect 186000 236898 186056 237134
rect 186292 236898 186348 237134
rect 186000 236866 186348 236898
rect 45234 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 45854 226894
rect 45234 226574 45854 226658
rect 45234 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 45854 226574
rect 45234 190894 45854 226338
rect 50952 219454 51300 219486
rect 50952 219218 51008 219454
rect 51244 219218 51300 219454
rect 50952 219134 51300 219218
rect 50952 218898 51008 219134
rect 51244 218898 51300 219134
rect 50952 218866 51300 218898
rect 185320 219454 185668 219486
rect 185320 219218 185376 219454
rect 185612 219218 185668 219454
rect 185320 219134 185668 219218
rect 185320 218898 185376 219134
rect 185612 218898 185668 219134
rect 185320 218866 185668 218898
rect 50272 201454 50620 201486
rect 50272 201218 50328 201454
rect 50564 201218 50620 201454
rect 50272 201134 50620 201218
rect 50272 200898 50328 201134
rect 50564 200898 50620 201134
rect 50272 200866 50620 200898
rect 186000 201454 186348 201486
rect 186000 201218 186056 201454
rect 186292 201218 186348 201454
rect 186000 201134 186348 201218
rect 186000 200898 186056 201134
rect 186292 200898 186348 201134
rect 186000 200866 186348 200898
rect 66056 199610 66116 200130
rect 67144 199610 67204 200130
rect 68232 199610 68292 200130
rect 69592 199610 69652 200130
rect 70544 199610 70604 200130
rect 66056 199550 66178 199610
rect 67144 199550 67282 199610
rect 68232 199550 68386 199610
rect 69592 199550 69674 199610
rect 45234 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 45854 190894
rect 45234 190574 45854 190658
rect 45234 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 45854 190574
rect 45234 154894 45854 190338
rect 45234 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 45854 154894
rect 45234 154574 45854 154658
rect 45234 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 45854 154574
rect 45234 118894 45854 154338
rect 45234 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 45854 118894
rect 45234 118574 45854 118658
rect 45234 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 45854 118574
rect 45234 82894 45854 118338
rect 45234 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 45854 82894
rect 45234 82574 45854 82658
rect 45234 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 45854 82574
rect 45234 46894 45854 82338
rect 45234 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 45854 46894
rect 45234 46574 45854 46658
rect 45234 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 45854 46574
rect 45234 10894 45854 46338
rect 45234 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 45854 10894
rect 45234 10574 45854 10658
rect 45234 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 45854 10574
rect 45234 -4186 45854 10338
rect 45234 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 45854 -4186
rect 45234 -4506 45854 -4422
rect 45234 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 45854 -4506
rect 45234 -5734 45854 -4742
rect 48954 194614 49574 198000
rect 48954 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 49574 194614
rect 48954 194294 49574 194378
rect 48954 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 49574 194294
rect 48954 158614 49574 194058
rect 48954 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 49574 158614
rect 48954 158294 49574 158378
rect 48954 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 49574 158294
rect 48954 122614 49574 158058
rect 48954 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 49574 122614
rect 48954 122294 49574 122378
rect 48954 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 49574 122294
rect 48954 86614 49574 122058
rect 48954 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 49574 86614
rect 48954 86294 49574 86378
rect 48954 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 49574 86294
rect 48954 50614 49574 86058
rect 48954 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 49574 50614
rect 48954 50294 49574 50378
rect 48954 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 49574 50294
rect 48954 14614 49574 50058
rect 48954 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 49574 14614
rect 48954 14294 49574 14378
rect 48954 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 49574 14294
rect 30954 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 31574 -7066
rect 30954 -7386 31574 -7302
rect 30954 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 31574 -7386
rect 30954 -7654 31574 -7622
rect 48954 -6106 49574 14058
rect 55794 165454 56414 198000
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -1306 56414 20898
rect 55794 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 56414 -1306
rect 55794 -1626 56414 -1542
rect 55794 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 56414 -1626
rect 55794 -1894 56414 -1862
rect 59514 169174 60134 198000
rect 59514 168938 59546 169174
rect 59782 168938 59866 169174
rect 60102 168938 60134 169174
rect 59514 168854 60134 168938
rect 59514 168618 59546 168854
rect 59782 168618 59866 168854
rect 60102 168618 60134 168854
rect 59514 133174 60134 168618
rect 59514 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 60134 133174
rect 59514 132854 60134 132938
rect 59514 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 60134 132854
rect 59514 97174 60134 132618
rect 59514 96938 59546 97174
rect 59782 96938 59866 97174
rect 60102 96938 60134 97174
rect 59514 96854 60134 96938
rect 59514 96618 59546 96854
rect 59782 96618 59866 96854
rect 60102 96618 60134 96854
rect 59514 61174 60134 96618
rect 59514 60938 59546 61174
rect 59782 60938 59866 61174
rect 60102 60938 60134 61174
rect 59514 60854 60134 60938
rect 59514 60618 59546 60854
rect 59782 60618 59866 60854
rect 60102 60618 60134 60854
rect 59514 25174 60134 60618
rect 59514 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 60134 25174
rect 59514 24854 60134 24938
rect 59514 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 60134 24854
rect 59514 -3226 60134 24618
rect 59514 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 60134 -3226
rect 59514 -3546 60134 -3462
rect 59514 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 60134 -3546
rect 59514 -3814 60134 -3782
rect 63234 172894 63854 198000
rect 66118 197437 66178 199550
rect 67222 198253 67282 199550
rect 67219 198252 67285 198253
rect 67219 198188 67220 198252
rect 67284 198188 67285 198252
rect 67219 198187 67285 198188
rect 66115 197436 66181 197437
rect 66115 197372 66116 197436
rect 66180 197372 66181 197436
rect 66115 197371 66181 197372
rect 63234 172658 63266 172894
rect 63502 172658 63586 172894
rect 63822 172658 63854 172894
rect 63234 172574 63854 172658
rect 63234 172338 63266 172574
rect 63502 172338 63586 172574
rect 63822 172338 63854 172574
rect 63234 136894 63854 172338
rect 63234 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 63854 136894
rect 63234 136574 63854 136658
rect 63234 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 63854 136574
rect 63234 100894 63854 136338
rect 63234 100658 63266 100894
rect 63502 100658 63586 100894
rect 63822 100658 63854 100894
rect 63234 100574 63854 100658
rect 63234 100338 63266 100574
rect 63502 100338 63586 100574
rect 63822 100338 63854 100574
rect 63234 64894 63854 100338
rect 63234 64658 63266 64894
rect 63502 64658 63586 64894
rect 63822 64658 63854 64894
rect 63234 64574 63854 64658
rect 63234 64338 63266 64574
rect 63502 64338 63586 64574
rect 63822 64338 63854 64574
rect 63234 28894 63854 64338
rect 63234 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 63854 28894
rect 63234 28574 63854 28658
rect 63234 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 63854 28574
rect 63234 -5146 63854 28338
rect 63234 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 63854 -5146
rect 63234 -5466 63854 -5382
rect 63234 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 63854 -5466
rect 63234 -5734 63854 -5702
rect 66954 176614 67574 198000
rect 68326 197437 68386 199550
rect 69614 197981 69674 199550
rect 70534 199550 70604 199610
rect 71768 199610 71828 200130
rect 73128 199610 73188 200130
rect 71768 199550 71882 199610
rect 70534 199477 70594 199550
rect 70531 199476 70597 199477
rect 70531 199412 70532 199476
rect 70596 199412 70597 199476
rect 70531 199411 70597 199412
rect 71822 198661 71882 199550
rect 73110 199550 73188 199610
rect 74214 200070 74276 200130
rect 71819 198660 71885 198661
rect 71819 198596 71820 198660
rect 71884 198596 71885 198660
rect 71819 198595 71885 198596
rect 73110 198389 73170 199550
rect 73107 198388 73173 198389
rect 73107 198324 73108 198388
rect 73172 198324 73173 198388
rect 73107 198323 73173 198324
rect 74214 198253 74274 200070
rect 75440 199610 75500 200130
rect 76528 199610 76588 200130
rect 77616 199610 77676 200130
rect 78296 199610 78356 200130
rect 75440 199550 75562 199610
rect 76528 199550 76666 199610
rect 77616 199550 77770 199610
rect 75502 198661 75562 199550
rect 76606 198661 76666 199550
rect 77710 199477 77770 199550
rect 78262 199550 78356 199610
rect 78704 199610 78764 200130
rect 80064 199610 80124 200130
rect 80744 199610 80804 200130
rect 81288 199610 81348 200130
rect 82376 199610 82436 200130
rect 83464 199610 83524 200130
rect 78704 199550 78874 199610
rect 80064 199550 80162 199610
rect 80744 199550 80898 199610
rect 81288 199550 81450 199610
rect 82376 199550 82554 199610
rect 77707 199476 77773 199477
rect 77707 199412 77708 199476
rect 77772 199412 77773 199476
rect 77707 199411 77773 199412
rect 75499 198660 75565 198661
rect 75499 198596 75500 198660
rect 75564 198596 75565 198660
rect 75499 198595 75565 198596
rect 76603 198660 76669 198661
rect 76603 198596 76604 198660
rect 76668 198596 76669 198660
rect 76603 198595 76669 198596
rect 74211 198252 74277 198253
rect 74211 198188 74212 198252
rect 74276 198188 74277 198252
rect 74211 198187 74277 198188
rect 69611 197980 69677 197981
rect 69611 197916 69612 197980
rect 69676 197916 69677 197980
rect 69611 197915 69677 197916
rect 68323 197436 68389 197437
rect 68323 197372 68324 197436
rect 68388 197372 68389 197436
rect 68323 197371 68389 197372
rect 66954 176378 66986 176614
rect 67222 176378 67306 176614
rect 67542 176378 67574 176614
rect 66954 176294 67574 176378
rect 66954 176058 66986 176294
rect 67222 176058 67306 176294
rect 67542 176058 67574 176294
rect 66954 140614 67574 176058
rect 66954 140378 66986 140614
rect 67222 140378 67306 140614
rect 67542 140378 67574 140614
rect 66954 140294 67574 140378
rect 66954 140058 66986 140294
rect 67222 140058 67306 140294
rect 67542 140058 67574 140294
rect 66954 104614 67574 140058
rect 66954 104378 66986 104614
rect 67222 104378 67306 104614
rect 67542 104378 67574 104614
rect 66954 104294 67574 104378
rect 66954 104058 66986 104294
rect 67222 104058 67306 104294
rect 67542 104058 67574 104294
rect 66954 68614 67574 104058
rect 66954 68378 66986 68614
rect 67222 68378 67306 68614
rect 67542 68378 67574 68614
rect 66954 68294 67574 68378
rect 66954 68058 66986 68294
rect 67222 68058 67306 68294
rect 67542 68058 67574 68294
rect 66954 32614 67574 68058
rect 66954 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 67574 32614
rect 66954 32294 67574 32378
rect 66954 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 67574 32294
rect 48954 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 49574 -6106
rect 48954 -6426 49574 -6342
rect 48954 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 49574 -6426
rect 48954 -7654 49574 -6662
rect 66954 -7066 67574 32058
rect 73794 183454 74414 198000
rect 73794 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 74414 183454
rect 73794 183134 74414 183218
rect 73794 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 74414 183134
rect 73794 147454 74414 182898
rect 73794 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 74414 147454
rect 73794 147134 74414 147218
rect 73794 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 74414 147134
rect 73794 111454 74414 146898
rect 73794 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 74414 111454
rect 73794 111134 74414 111218
rect 73794 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 74414 111134
rect 73794 75454 74414 110898
rect 73794 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 74414 75454
rect 73794 75134 74414 75218
rect 73794 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 74414 75134
rect 73794 39454 74414 74898
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -1894 74414 -902
rect 77514 187174 78134 198000
rect 78262 197437 78322 199550
rect 78814 199477 78874 199550
rect 78811 199476 78877 199477
rect 78811 199412 78812 199476
rect 78876 199412 78877 199476
rect 78811 199411 78877 199412
rect 80102 198661 80162 199550
rect 80099 198660 80165 198661
rect 80099 198596 80100 198660
rect 80164 198596 80165 198660
rect 80099 198595 80165 198596
rect 80838 197437 80898 199550
rect 81390 198661 81450 199550
rect 82494 198661 82554 199550
rect 83414 199550 83524 199610
rect 83598 200070 83660 200130
rect 81387 198660 81453 198661
rect 81387 198596 81388 198660
rect 81452 198596 81453 198660
rect 81387 198595 81453 198596
rect 82491 198660 82557 198661
rect 82491 198596 82492 198660
rect 82556 198596 82557 198660
rect 82491 198595 82557 198596
rect 83414 198389 83474 199550
rect 83411 198388 83477 198389
rect 83411 198324 83412 198388
rect 83476 198324 83477 198388
rect 83411 198323 83477 198324
rect 83598 198253 83658 200070
rect 84552 199610 84612 200130
rect 85912 199610 85972 200130
rect 84518 199550 84612 199610
rect 85806 199550 85972 199610
rect 86048 199610 86108 200130
rect 87000 199610 87060 200130
rect 88088 199610 88148 200130
rect 88496 199610 88556 200130
rect 89448 199610 89508 200130
rect 90672 199610 90732 200130
rect 91080 199610 91140 200130
rect 91760 199610 91820 200130
rect 92848 199610 92908 200130
rect 93528 200070 93594 200130
rect 86048 199550 86234 199610
rect 87000 199550 87154 199610
rect 88088 199550 88258 199610
rect 88496 199550 88626 199610
rect 89448 199550 89546 199610
rect 90672 199550 90834 199610
rect 91080 199550 91202 199610
rect 84518 198661 84578 199550
rect 84515 198660 84581 198661
rect 84515 198596 84516 198660
rect 84580 198596 84581 198660
rect 84515 198595 84581 198596
rect 85806 198525 85866 199550
rect 86174 198661 86234 199550
rect 87094 198661 87154 199550
rect 86171 198660 86237 198661
rect 86171 198596 86172 198660
rect 86236 198596 86237 198660
rect 86171 198595 86237 198596
rect 87091 198660 87157 198661
rect 87091 198596 87092 198660
rect 87156 198596 87157 198660
rect 87091 198595 87157 198596
rect 88198 198525 88258 199550
rect 88566 199477 88626 199550
rect 88563 199476 88629 199477
rect 88563 199412 88564 199476
rect 88628 199412 88629 199476
rect 88563 199411 88629 199412
rect 89486 198525 89546 199550
rect 90774 198525 90834 199550
rect 91142 199477 91202 199550
rect 91510 199550 91820 199610
rect 92798 199550 92908 199610
rect 91139 199476 91205 199477
rect 91139 199412 91140 199476
rect 91204 199412 91205 199476
rect 91139 199411 91205 199412
rect 85803 198524 85869 198525
rect 85803 198460 85804 198524
rect 85868 198460 85869 198524
rect 85803 198459 85869 198460
rect 88195 198524 88261 198525
rect 88195 198460 88196 198524
rect 88260 198460 88261 198524
rect 88195 198459 88261 198460
rect 89483 198524 89549 198525
rect 89483 198460 89484 198524
rect 89548 198460 89549 198524
rect 89483 198459 89549 198460
rect 90771 198524 90837 198525
rect 90771 198460 90772 198524
rect 90836 198460 90837 198524
rect 90771 198459 90837 198460
rect 83595 198252 83661 198253
rect 83595 198188 83596 198252
rect 83660 198188 83661 198252
rect 83595 198187 83661 198188
rect 78259 197436 78325 197437
rect 78259 197372 78260 197436
rect 78324 197372 78325 197436
rect 78259 197371 78325 197372
rect 80835 197436 80901 197437
rect 80835 197372 80836 197436
rect 80900 197372 80901 197436
rect 80835 197371 80901 197372
rect 77514 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 78134 187174
rect 77514 186854 78134 186938
rect 77514 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 78134 186854
rect 77514 151174 78134 186618
rect 77514 150938 77546 151174
rect 77782 150938 77866 151174
rect 78102 150938 78134 151174
rect 77514 150854 78134 150938
rect 77514 150618 77546 150854
rect 77782 150618 77866 150854
rect 78102 150618 78134 150854
rect 77514 115174 78134 150618
rect 77514 114938 77546 115174
rect 77782 114938 77866 115174
rect 78102 114938 78134 115174
rect 77514 114854 78134 114938
rect 77514 114618 77546 114854
rect 77782 114618 77866 114854
rect 78102 114618 78134 114854
rect 77514 79174 78134 114618
rect 77514 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 78134 79174
rect 77514 78854 78134 78938
rect 77514 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 78134 78854
rect 77514 43174 78134 78618
rect 77514 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 78134 43174
rect 77514 42854 78134 42938
rect 77514 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 78134 42854
rect 77514 7174 78134 42618
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -2266 78134 6618
rect 77514 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 78134 -2266
rect 77514 -2586 78134 -2502
rect 77514 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 78134 -2586
rect 77514 -3814 78134 -2822
rect 81234 190894 81854 198000
rect 81234 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 81854 190894
rect 81234 190574 81854 190658
rect 81234 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 81854 190574
rect 81234 154894 81854 190338
rect 81234 154658 81266 154894
rect 81502 154658 81586 154894
rect 81822 154658 81854 154894
rect 81234 154574 81854 154658
rect 81234 154338 81266 154574
rect 81502 154338 81586 154574
rect 81822 154338 81854 154574
rect 81234 118894 81854 154338
rect 81234 118658 81266 118894
rect 81502 118658 81586 118894
rect 81822 118658 81854 118894
rect 81234 118574 81854 118658
rect 81234 118338 81266 118574
rect 81502 118338 81586 118574
rect 81822 118338 81854 118574
rect 81234 82894 81854 118338
rect 81234 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 81854 82894
rect 81234 82574 81854 82658
rect 81234 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 81854 82574
rect 81234 46894 81854 82338
rect 81234 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 81854 46894
rect 81234 46574 81854 46658
rect 81234 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 81854 46574
rect 81234 10894 81854 46338
rect 81234 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 81854 10894
rect 81234 10574 81854 10658
rect 81234 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 81854 10574
rect 81234 -4186 81854 10338
rect 81234 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 81854 -4186
rect 81234 -4506 81854 -4422
rect 81234 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 81854 -4506
rect 81234 -5734 81854 -4742
rect 84954 194614 85574 198000
rect 91510 197573 91570 199550
rect 92798 198661 92858 199550
rect 93534 198661 93594 200070
rect 93936 199610 93996 200130
rect 93902 199550 93996 199610
rect 95296 199610 95356 200130
rect 95976 199610 96036 200130
rect 95296 199550 95434 199610
rect 92795 198660 92861 198661
rect 92795 198596 92796 198660
rect 92860 198596 92861 198660
rect 92795 198595 92861 198596
rect 93531 198660 93597 198661
rect 93531 198596 93532 198660
rect 93596 198596 93597 198660
rect 93531 198595 93597 198596
rect 93902 198253 93962 199550
rect 93899 198252 93965 198253
rect 93899 198188 93900 198252
rect 93964 198188 93965 198252
rect 93899 198187 93965 198188
rect 95374 198117 95434 199550
rect 95926 199550 96036 199610
rect 96384 199610 96444 200130
rect 97608 199610 97668 200130
rect 96384 199550 96538 199610
rect 95926 198661 95986 199550
rect 96478 198933 96538 199550
rect 97582 199550 97668 199610
rect 98288 199610 98348 200130
rect 98696 199610 98756 200130
rect 99784 200070 99850 200130
rect 98288 199550 98378 199610
rect 96475 198932 96541 198933
rect 96475 198868 96476 198932
rect 96540 198868 96541 198932
rect 96475 198867 96541 198868
rect 97582 198661 97642 199550
rect 95923 198660 95989 198661
rect 95923 198596 95924 198660
rect 95988 198596 95989 198660
rect 95923 198595 95989 198596
rect 97579 198660 97645 198661
rect 97579 198596 97580 198660
rect 97644 198596 97645 198660
rect 97579 198595 97645 198596
rect 98318 198525 98378 199550
rect 98686 199550 98756 199610
rect 98686 199069 98746 199550
rect 98683 199068 98749 199069
rect 98683 199004 98684 199068
rect 98748 199004 98749 199068
rect 98683 199003 98749 199004
rect 99790 198525 99850 200070
rect 101008 199610 101068 200130
rect 100894 199550 101068 199610
rect 101144 199610 101204 200130
rect 102232 199610 102292 200130
rect 103320 199610 103380 200130
rect 101144 199550 101322 199610
rect 100894 198525 100954 199550
rect 98315 198524 98381 198525
rect 98315 198460 98316 198524
rect 98380 198460 98381 198524
rect 98315 198459 98381 198460
rect 99787 198524 99853 198525
rect 99787 198460 99788 198524
rect 99852 198460 99853 198524
rect 99787 198459 99853 198460
rect 100891 198524 100957 198525
rect 100891 198460 100892 198524
rect 100956 198460 100957 198524
rect 100891 198459 100957 198460
rect 95371 198116 95437 198117
rect 95371 198052 95372 198116
rect 95436 198052 95437 198116
rect 95371 198051 95437 198052
rect 91507 197572 91573 197573
rect 91507 197508 91508 197572
rect 91572 197508 91573 197572
rect 91507 197507 91573 197508
rect 84954 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 85574 194614
rect 84954 194294 85574 194378
rect 84954 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 85574 194294
rect 84954 158614 85574 194058
rect 84954 158378 84986 158614
rect 85222 158378 85306 158614
rect 85542 158378 85574 158614
rect 84954 158294 85574 158378
rect 84954 158058 84986 158294
rect 85222 158058 85306 158294
rect 85542 158058 85574 158294
rect 84954 122614 85574 158058
rect 84954 122378 84986 122614
rect 85222 122378 85306 122614
rect 85542 122378 85574 122614
rect 84954 122294 85574 122378
rect 84954 122058 84986 122294
rect 85222 122058 85306 122294
rect 85542 122058 85574 122294
rect 84954 86614 85574 122058
rect 84954 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 85574 86614
rect 84954 86294 85574 86378
rect 84954 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 85574 86294
rect 84954 50614 85574 86058
rect 84954 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 85574 50614
rect 84954 50294 85574 50378
rect 84954 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 85574 50294
rect 84954 14614 85574 50058
rect 84954 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 85574 14614
rect 84954 14294 85574 14378
rect 84954 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 85574 14294
rect 66954 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 67574 -7066
rect 66954 -7386 67574 -7302
rect 66954 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 67574 -7386
rect 66954 -7654 67574 -7622
rect 84954 -6106 85574 14058
rect 91794 165454 92414 198000
rect 91794 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 92414 165454
rect 91794 165134 92414 165218
rect 91794 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 92414 165134
rect 91794 129454 92414 164898
rect 91794 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 92414 129454
rect 91794 129134 92414 129218
rect 91794 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 92414 129134
rect 91794 93454 92414 128898
rect 91794 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 92414 93454
rect 91794 93134 92414 93218
rect 91794 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 92414 93134
rect 91794 57454 92414 92898
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -1306 92414 20898
rect 91794 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 92414 -1306
rect 91794 -1626 92414 -1542
rect 91794 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 92414 -1626
rect 91794 -1894 92414 -1862
rect 95514 169174 96134 198000
rect 95514 168938 95546 169174
rect 95782 168938 95866 169174
rect 96102 168938 96134 169174
rect 95514 168854 96134 168938
rect 95514 168618 95546 168854
rect 95782 168618 95866 168854
rect 96102 168618 96134 168854
rect 95514 133174 96134 168618
rect 95514 132938 95546 133174
rect 95782 132938 95866 133174
rect 96102 132938 96134 133174
rect 95514 132854 96134 132938
rect 95514 132618 95546 132854
rect 95782 132618 95866 132854
rect 96102 132618 96134 132854
rect 95514 97174 96134 132618
rect 95514 96938 95546 97174
rect 95782 96938 95866 97174
rect 96102 96938 96134 97174
rect 95514 96854 96134 96938
rect 95514 96618 95546 96854
rect 95782 96618 95866 96854
rect 96102 96618 96134 96854
rect 95514 61174 96134 96618
rect 95514 60938 95546 61174
rect 95782 60938 95866 61174
rect 96102 60938 96134 61174
rect 95514 60854 96134 60938
rect 95514 60618 95546 60854
rect 95782 60618 95866 60854
rect 96102 60618 96134 60854
rect 95514 25174 96134 60618
rect 95514 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 96134 25174
rect 95514 24854 96134 24938
rect 95514 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 96134 24854
rect 95514 -3226 96134 24618
rect 95514 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 96134 -3226
rect 95514 -3546 96134 -3462
rect 95514 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 96134 -3546
rect 95514 -3814 96134 -3782
rect 99234 172894 99854 198000
rect 101262 197165 101322 199550
rect 102182 199550 102292 199610
rect 103286 199550 103380 199610
rect 103592 199610 103652 200130
rect 104408 199610 104468 200130
rect 103592 199550 103714 199610
rect 102182 198525 102242 199550
rect 103286 198525 103346 199550
rect 103654 199477 103714 199550
rect 104390 199550 104468 199610
rect 105768 199610 105828 200130
rect 106040 200070 106106 200130
rect 105768 199550 105922 199610
rect 103651 199476 103717 199477
rect 103651 199412 103652 199476
rect 103716 199412 103717 199476
rect 103651 199411 103717 199412
rect 104390 198661 104450 199550
rect 105862 198661 105922 199550
rect 106046 198661 106106 200070
rect 106992 199610 107052 200130
rect 108080 199610 108140 200130
rect 108488 199610 108548 200130
rect 109168 200070 109234 200130
rect 106966 199550 107052 199610
rect 108070 199550 108140 199610
rect 108438 199550 108548 199610
rect 104387 198660 104453 198661
rect 104387 198596 104388 198660
rect 104452 198596 104453 198660
rect 104387 198595 104453 198596
rect 105859 198660 105925 198661
rect 105859 198596 105860 198660
rect 105924 198596 105925 198660
rect 105859 198595 105925 198596
rect 106043 198660 106109 198661
rect 106043 198596 106044 198660
rect 106108 198596 106109 198660
rect 106043 198595 106109 198596
rect 102179 198524 102245 198525
rect 102179 198460 102180 198524
rect 102244 198460 102245 198524
rect 102179 198459 102245 198460
rect 103283 198524 103349 198525
rect 103283 198460 103284 198524
rect 103348 198460 103349 198524
rect 103283 198459 103349 198460
rect 101259 197164 101325 197165
rect 101259 197100 101260 197164
rect 101324 197100 101325 197164
rect 101259 197099 101325 197100
rect 99234 172658 99266 172894
rect 99502 172658 99586 172894
rect 99822 172658 99854 172894
rect 99234 172574 99854 172658
rect 99234 172338 99266 172574
rect 99502 172338 99586 172574
rect 99822 172338 99854 172574
rect 99234 136894 99854 172338
rect 99234 136658 99266 136894
rect 99502 136658 99586 136894
rect 99822 136658 99854 136894
rect 99234 136574 99854 136658
rect 99234 136338 99266 136574
rect 99502 136338 99586 136574
rect 99822 136338 99854 136574
rect 99234 100894 99854 136338
rect 99234 100658 99266 100894
rect 99502 100658 99586 100894
rect 99822 100658 99854 100894
rect 99234 100574 99854 100658
rect 99234 100338 99266 100574
rect 99502 100338 99586 100574
rect 99822 100338 99854 100574
rect 99234 64894 99854 100338
rect 99234 64658 99266 64894
rect 99502 64658 99586 64894
rect 99822 64658 99854 64894
rect 99234 64574 99854 64658
rect 99234 64338 99266 64574
rect 99502 64338 99586 64574
rect 99822 64338 99854 64574
rect 99234 28894 99854 64338
rect 99234 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 99854 28894
rect 99234 28574 99854 28658
rect 99234 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 99854 28574
rect 99234 -5146 99854 28338
rect 99234 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 99854 -5146
rect 99234 -5466 99854 -5382
rect 99234 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 99854 -5466
rect 99234 -5734 99854 -5702
rect 102954 176614 103574 198000
rect 106966 197981 107026 199550
rect 108070 197981 108130 199550
rect 108438 198661 108498 199550
rect 108435 198660 108501 198661
rect 108435 198596 108436 198660
rect 108500 198596 108501 198660
rect 108435 198595 108501 198596
rect 109174 197981 109234 200070
rect 110936 199610 110996 200130
rect 113520 199610 113580 200130
rect 115968 199610 116028 200130
rect 118280 199610 118340 200130
rect 121000 199610 121060 200130
rect 110936 199550 111074 199610
rect 113520 199550 113650 199610
rect 115968 199550 116042 199610
rect 118280 199550 118434 199610
rect 111014 199477 111074 199550
rect 111011 199476 111077 199477
rect 111011 199412 111012 199476
rect 111076 199412 111077 199476
rect 111011 199411 111077 199412
rect 113590 198661 113650 199550
rect 115982 198661 116042 199550
rect 118374 198661 118434 199550
rect 120950 199550 121060 199610
rect 123448 199610 123508 200130
rect 125896 199610 125956 200130
rect 128480 199610 128540 200130
rect 130928 199610 130988 200130
rect 133512 199610 133572 200130
rect 123448 199550 123586 199610
rect 125896 199550 125978 199610
rect 128480 199550 128554 199610
rect 120950 198661 121010 199550
rect 123526 198661 123586 199550
rect 125918 198661 125978 199550
rect 128494 198661 128554 199550
rect 130886 199550 130988 199610
rect 133462 199550 133572 199610
rect 135960 199610 136020 200130
rect 138544 199610 138604 200130
rect 140992 199610 141052 200130
rect 143440 199610 143500 200130
rect 135960 199550 136098 199610
rect 138544 199550 138674 199610
rect 140992 199550 141066 199610
rect 113587 198660 113653 198661
rect 113587 198596 113588 198660
rect 113652 198596 113653 198660
rect 113587 198595 113653 198596
rect 115979 198660 116045 198661
rect 115979 198596 115980 198660
rect 116044 198596 116045 198660
rect 115979 198595 116045 198596
rect 118371 198660 118437 198661
rect 118371 198596 118372 198660
rect 118436 198596 118437 198660
rect 118371 198595 118437 198596
rect 120947 198660 121013 198661
rect 120947 198596 120948 198660
rect 121012 198596 121013 198660
rect 120947 198595 121013 198596
rect 123523 198660 123589 198661
rect 123523 198596 123524 198660
rect 123588 198596 123589 198660
rect 123523 198595 123589 198596
rect 125915 198660 125981 198661
rect 125915 198596 125916 198660
rect 125980 198596 125981 198660
rect 125915 198595 125981 198596
rect 128491 198660 128557 198661
rect 128491 198596 128492 198660
rect 128556 198596 128557 198660
rect 128491 198595 128557 198596
rect 106963 197980 107029 197981
rect 106963 197916 106964 197980
rect 107028 197916 107029 197980
rect 106963 197915 107029 197916
rect 108067 197980 108133 197981
rect 108067 197916 108068 197980
rect 108132 197916 108133 197980
rect 108067 197915 108133 197916
rect 109171 197980 109237 197981
rect 109171 197916 109172 197980
rect 109236 197916 109237 197980
rect 109171 197915 109237 197916
rect 102954 176378 102986 176614
rect 103222 176378 103306 176614
rect 103542 176378 103574 176614
rect 102954 176294 103574 176378
rect 102954 176058 102986 176294
rect 103222 176058 103306 176294
rect 103542 176058 103574 176294
rect 102954 140614 103574 176058
rect 102954 140378 102986 140614
rect 103222 140378 103306 140614
rect 103542 140378 103574 140614
rect 102954 140294 103574 140378
rect 102954 140058 102986 140294
rect 103222 140058 103306 140294
rect 103542 140058 103574 140294
rect 102954 104614 103574 140058
rect 102954 104378 102986 104614
rect 103222 104378 103306 104614
rect 103542 104378 103574 104614
rect 102954 104294 103574 104378
rect 102954 104058 102986 104294
rect 103222 104058 103306 104294
rect 103542 104058 103574 104294
rect 102954 68614 103574 104058
rect 102954 68378 102986 68614
rect 103222 68378 103306 68614
rect 103542 68378 103574 68614
rect 102954 68294 103574 68378
rect 102954 68058 102986 68294
rect 103222 68058 103306 68294
rect 103542 68058 103574 68294
rect 102954 32614 103574 68058
rect 102954 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 103574 32614
rect 102954 32294 103574 32378
rect 102954 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 103574 32294
rect 84954 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 85574 -6106
rect 84954 -6426 85574 -6342
rect 84954 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 85574 -6426
rect 84954 -7654 85574 -6662
rect 102954 -7066 103574 32058
rect 109794 183454 110414 198000
rect 109794 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 110414 183454
rect 109794 183134 110414 183218
rect 109794 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 110414 183134
rect 109794 147454 110414 182898
rect 109794 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 110414 147454
rect 109794 147134 110414 147218
rect 109794 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 110414 147134
rect 109794 111454 110414 146898
rect 109794 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 110414 111454
rect 109794 111134 110414 111218
rect 109794 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 110414 111134
rect 109794 75454 110414 110898
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 109794 39454 110414 74898
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -1894 110414 -902
rect 113514 187174 114134 198000
rect 113514 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 114134 187174
rect 113514 186854 114134 186938
rect 113514 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 114134 186854
rect 113514 151174 114134 186618
rect 113514 150938 113546 151174
rect 113782 150938 113866 151174
rect 114102 150938 114134 151174
rect 113514 150854 114134 150938
rect 113514 150618 113546 150854
rect 113782 150618 113866 150854
rect 114102 150618 114134 150854
rect 113514 115174 114134 150618
rect 113514 114938 113546 115174
rect 113782 114938 113866 115174
rect 114102 114938 114134 115174
rect 113514 114854 114134 114938
rect 113514 114618 113546 114854
rect 113782 114618 113866 114854
rect 114102 114618 114134 114854
rect 113514 79174 114134 114618
rect 113514 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 114134 79174
rect 113514 78854 114134 78938
rect 113514 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 114134 78854
rect 113514 43174 114134 78618
rect 113514 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 114134 43174
rect 113514 42854 114134 42938
rect 113514 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 114134 42854
rect 113514 7174 114134 42618
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 113514 -2266 114134 6618
rect 113514 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 114134 -2266
rect 113514 -2586 114134 -2502
rect 113514 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 114134 -2586
rect 113514 -3814 114134 -2822
rect 117234 190894 117854 198000
rect 117234 190658 117266 190894
rect 117502 190658 117586 190894
rect 117822 190658 117854 190894
rect 117234 190574 117854 190658
rect 117234 190338 117266 190574
rect 117502 190338 117586 190574
rect 117822 190338 117854 190574
rect 117234 154894 117854 190338
rect 117234 154658 117266 154894
rect 117502 154658 117586 154894
rect 117822 154658 117854 154894
rect 117234 154574 117854 154658
rect 117234 154338 117266 154574
rect 117502 154338 117586 154574
rect 117822 154338 117854 154574
rect 117234 118894 117854 154338
rect 117234 118658 117266 118894
rect 117502 118658 117586 118894
rect 117822 118658 117854 118894
rect 117234 118574 117854 118658
rect 117234 118338 117266 118574
rect 117502 118338 117586 118574
rect 117822 118338 117854 118574
rect 117234 82894 117854 118338
rect 117234 82658 117266 82894
rect 117502 82658 117586 82894
rect 117822 82658 117854 82894
rect 117234 82574 117854 82658
rect 117234 82338 117266 82574
rect 117502 82338 117586 82574
rect 117822 82338 117854 82574
rect 117234 46894 117854 82338
rect 117234 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 117854 46894
rect 117234 46574 117854 46658
rect 117234 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 117854 46574
rect 117234 10894 117854 46338
rect 117234 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 117854 10894
rect 117234 10574 117854 10658
rect 117234 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 117854 10574
rect 117234 -4186 117854 10338
rect 117234 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 117854 -4186
rect 117234 -4506 117854 -4422
rect 117234 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 117854 -4506
rect 117234 -5734 117854 -4742
rect 120954 194614 121574 198000
rect 120954 194378 120986 194614
rect 121222 194378 121306 194614
rect 121542 194378 121574 194614
rect 120954 194294 121574 194378
rect 120954 194058 120986 194294
rect 121222 194058 121306 194294
rect 121542 194058 121574 194294
rect 120954 158614 121574 194058
rect 120954 158378 120986 158614
rect 121222 158378 121306 158614
rect 121542 158378 121574 158614
rect 120954 158294 121574 158378
rect 120954 158058 120986 158294
rect 121222 158058 121306 158294
rect 121542 158058 121574 158294
rect 120954 122614 121574 158058
rect 120954 122378 120986 122614
rect 121222 122378 121306 122614
rect 121542 122378 121574 122614
rect 120954 122294 121574 122378
rect 120954 122058 120986 122294
rect 121222 122058 121306 122294
rect 121542 122058 121574 122294
rect 120954 86614 121574 122058
rect 120954 86378 120986 86614
rect 121222 86378 121306 86614
rect 121542 86378 121574 86614
rect 120954 86294 121574 86378
rect 120954 86058 120986 86294
rect 121222 86058 121306 86294
rect 121542 86058 121574 86294
rect 120954 50614 121574 86058
rect 120954 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 121574 50614
rect 120954 50294 121574 50378
rect 120954 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 121574 50294
rect 120954 14614 121574 50058
rect 120954 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 121574 14614
rect 120954 14294 121574 14378
rect 120954 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 121574 14294
rect 102954 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 103574 -7066
rect 102954 -7386 103574 -7302
rect 102954 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 103574 -7386
rect 102954 -7654 103574 -7622
rect 120954 -6106 121574 14058
rect 127794 165454 128414 198000
rect 130886 197981 130946 199550
rect 130883 197980 130949 197981
rect 130883 197916 130884 197980
rect 130948 197916 130949 197980
rect 130883 197915 130949 197916
rect 127794 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 128414 165454
rect 127794 165134 128414 165218
rect 127794 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 128414 165134
rect 127794 129454 128414 164898
rect 127794 129218 127826 129454
rect 128062 129218 128146 129454
rect 128382 129218 128414 129454
rect 127794 129134 128414 129218
rect 127794 128898 127826 129134
rect 128062 128898 128146 129134
rect 128382 128898 128414 129134
rect 127794 93454 128414 128898
rect 127794 93218 127826 93454
rect 128062 93218 128146 93454
rect 128382 93218 128414 93454
rect 127794 93134 128414 93218
rect 127794 92898 127826 93134
rect 128062 92898 128146 93134
rect 128382 92898 128414 93134
rect 127794 57454 128414 92898
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -1306 128414 20898
rect 127794 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 128414 -1306
rect 127794 -1626 128414 -1542
rect 127794 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 128414 -1626
rect 127794 -1894 128414 -1862
rect 131514 169174 132134 198000
rect 133462 197709 133522 199550
rect 136038 198797 136098 199550
rect 136035 198796 136101 198797
rect 136035 198732 136036 198796
rect 136100 198732 136101 198796
rect 136035 198731 136101 198732
rect 133459 197708 133525 197709
rect 133459 197644 133460 197708
rect 133524 197644 133525 197708
rect 133459 197643 133525 197644
rect 131514 168938 131546 169174
rect 131782 168938 131866 169174
rect 132102 168938 132134 169174
rect 131514 168854 132134 168938
rect 131514 168618 131546 168854
rect 131782 168618 131866 168854
rect 132102 168618 132134 168854
rect 131514 133174 132134 168618
rect 131514 132938 131546 133174
rect 131782 132938 131866 133174
rect 132102 132938 132134 133174
rect 131514 132854 132134 132938
rect 131514 132618 131546 132854
rect 131782 132618 131866 132854
rect 132102 132618 132134 132854
rect 131514 97174 132134 132618
rect 131514 96938 131546 97174
rect 131782 96938 131866 97174
rect 132102 96938 132134 97174
rect 131514 96854 132134 96938
rect 131514 96618 131546 96854
rect 131782 96618 131866 96854
rect 132102 96618 132134 96854
rect 131514 61174 132134 96618
rect 131514 60938 131546 61174
rect 131782 60938 131866 61174
rect 132102 60938 132134 61174
rect 131514 60854 132134 60938
rect 131514 60618 131546 60854
rect 131782 60618 131866 60854
rect 132102 60618 132134 60854
rect 131514 25174 132134 60618
rect 131514 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 132134 25174
rect 131514 24854 132134 24938
rect 131514 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 132134 24854
rect 131514 -3226 132134 24618
rect 131514 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 132134 -3226
rect 131514 -3546 132134 -3462
rect 131514 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 132134 -3546
rect 131514 -3814 132134 -3782
rect 135234 172894 135854 198000
rect 138614 197845 138674 199550
rect 138611 197844 138677 197845
rect 138611 197780 138612 197844
rect 138676 197780 138677 197844
rect 138611 197779 138677 197780
rect 135234 172658 135266 172894
rect 135502 172658 135586 172894
rect 135822 172658 135854 172894
rect 135234 172574 135854 172658
rect 135234 172338 135266 172574
rect 135502 172338 135586 172574
rect 135822 172338 135854 172574
rect 135234 136894 135854 172338
rect 135234 136658 135266 136894
rect 135502 136658 135586 136894
rect 135822 136658 135854 136894
rect 135234 136574 135854 136658
rect 135234 136338 135266 136574
rect 135502 136338 135586 136574
rect 135822 136338 135854 136574
rect 135234 100894 135854 136338
rect 135234 100658 135266 100894
rect 135502 100658 135586 100894
rect 135822 100658 135854 100894
rect 135234 100574 135854 100658
rect 135234 100338 135266 100574
rect 135502 100338 135586 100574
rect 135822 100338 135854 100574
rect 135234 64894 135854 100338
rect 135234 64658 135266 64894
rect 135502 64658 135586 64894
rect 135822 64658 135854 64894
rect 135234 64574 135854 64658
rect 135234 64338 135266 64574
rect 135502 64338 135586 64574
rect 135822 64338 135854 64574
rect 135234 28894 135854 64338
rect 135234 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 135854 28894
rect 135234 28574 135854 28658
rect 135234 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 135854 28574
rect 135234 -5146 135854 28338
rect 135234 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 135854 -5146
rect 135234 -5466 135854 -5382
rect 135234 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 135854 -5466
rect 135234 -5734 135854 -5702
rect 138954 176614 139574 198000
rect 141006 197845 141066 199550
rect 143398 199550 143500 199610
rect 145888 199610 145948 200130
rect 148472 199610 148532 200130
rect 150920 199610 150980 200130
rect 153368 199610 153428 200130
rect 155952 199610 156012 200130
rect 173224 199610 173284 200130
rect 145888 199550 146034 199610
rect 148472 199550 148610 199610
rect 150920 199550 151002 199610
rect 143398 197845 143458 199550
rect 145974 198661 146034 199550
rect 145971 198660 146037 198661
rect 145971 198596 145972 198660
rect 146036 198596 146037 198660
rect 145971 198595 146037 198596
rect 141003 197844 141069 197845
rect 141003 197780 141004 197844
rect 141068 197780 141069 197844
rect 141003 197779 141069 197780
rect 143395 197844 143461 197845
rect 143395 197780 143396 197844
rect 143460 197780 143461 197844
rect 143395 197779 143461 197780
rect 138954 176378 138986 176614
rect 139222 176378 139306 176614
rect 139542 176378 139574 176614
rect 138954 176294 139574 176378
rect 138954 176058 138986 176294
rect 139222 176058 139306 176294
rect 139542 176058 139574 176294
rect 138954 140614 139574 176058
rect 138954 140378 138986 140614
rect 139222 140378 139306 140614
rect 139542 140378 139574 140614
rect 138954 140294 139574 140378
rect 138954 140058 138986 140294
rect 139222 140058 139306 140294
rect 139542 140058 139574 140294
rect 138954 104614 139574 140058
rect 138954 104378 138986 104614
rect 139222 104378 139306 104614
rect 139542 104378 139574 104614
rect 138954 104294 139574 104378
rect 138954 104058 138986 104294
rect 139222 104058 139306 104294
rect 139542 104058 139574 104294
rect 138954 68614 139574 104058
rect 138954 68378 138986 68614
rect 139222 68378 139306 68614
rect 139542 68378 139574 68614
rect 138954 68294 139574 68378
rect 138954 68058 138986 68294
rect 139222 68058 139306 68294
rect 139542 68058 139574 68294
rect 138954 32614 139574 68058
rect 138954 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 139574 32614
rect 138954 32294 139574 32378
rect 138954 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 139574 32294
rect 120954 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 121574 -6106
rect 120954 -6426 121574 -6342
rect 120954 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 121574 -6426
rect 120954 -7654 121574 -6662
rect 138954 -7066 139574 32058
rect 145794 183454 146414 198000
rect 148550 197709 148610 199550
rect 148547 197708 148613 197709
rect 148547 197644 148548 197708
rect 148612 197644 148613 197708
rect 148547 197643 148613 197644
rect 145794 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 146414 183454
rect 145794 183134 146414 183218
rect 145794 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 146414 183134
rect 145794 147454 146414 182898
rect 145794 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 146414 147454
rect 145794 147134 146414 147218
rect 145794 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 146414 147134
rect 145794 111454 146414 146898
rect 145794 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 146414 111454
rect 145794 111134 146414 111218
rect 145794 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 146414 111134
rect 145794 75454 146414 110898
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 145794 39454 146414 74898
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -1894 146414 -902
rect 149514 187174 150134 198000
rect 150942 197709 151002 199550
rect 153334 199550 153428 199610
rect 155910 199550 156012 199610
rect 173206 199550 173284 199610
rect 173360 199610 173420 200130
rect 173360 199550 173450 199610
rect 153334 198661 153394 199550
rect 153331 198660 153397 198661
rect 153331 198596 153332 198660
rect 153396 198596 153397 198660
rect 153331 198595 153397 198596
rect 150939 197708 151005 197709
rect 150939 197644 150940 197708
rect 151004 197644 151005 197708
rect 150939 197643 151005 197644
rect 149514 186938 149546 187174
rect 149782 186938 149866 187174
rect 150102 186938 150134 187174
rect 149514 186854 150134 186938
rect 149514 186618 149546 186854
rect 149782 186618 149866 186854
rect 150102 186618 150134 186854
rect 149514 151174 150134 186618
rect 149514 150938 149546 151174
rect 149782 150938 149866 151174
rect 150102 150938 150134 151174
rect 149514 150854 150134 150938
rect 149514 150618 149546 150854
rect 149782 150618 149866 150854
rect 150102 150618 150134 150854
rect 149514 115174 150134 150618
rect 149514 114938 149546 115174
rect 149782 114938 149866 115174
rect 150102 114938 150134 115174
rect 149514 114854 150134 114938
rect 149514 114618 149546 114854
rect 149782 114618 149866 114854
rect 150102 114618 150134 114854
rect 149514 79174 150134 114618
rect 149514 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 150134 79174
rect 149514 78854 150134 78938
rect 149514 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 150134 78854
rect 149514 43174 150134 78618
rect 149514 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 150134 43174
rect 149514 42854 150134 42938
rect 149514 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 150134 42854
rect 149514 7174 150134 42618
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -2266 150134 6618
rect 149514 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 150134 -2266
rect 149514 -2586 150134 -2502
rect 149514 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 150134 -2586
rect 149514 -3814 150134 -2822
rect 153234 190894 153854 198000
rect 155910 197437 155970 199550
rect 155907 197436 155973 197437
rect 155907 197372 155908 197436
rect 155972 197372 155973 197436
rect 155907 197371 155973 197372
rect 153234 190658 153266 190894
rect 153502 190658 153586 190894
rect 153822 190658 153854 190894
rect 153234 190574 153854 190658
rect 153234 190338 153266 190574
rect 153502 190338 153586 190574
rect 153822 190338 153854 190574
rect 153234 154894 153854 190338
rect 153234 154658 153266 154894
rect 153502 154658 153586 154894
rect 153822 154658 153854 154894
rect 153234 154574 153854 154658
rect 153234 154338 153266 154574
rect 153502 154338 153586 154574
rect 153822 154338 153854 154574
rect 153234 118894 153854 154338
rect 153234 118658 153266 118894
rect 153502 118658 153586 118894
rect 153822 118658 153854 118894
rect 153234 118574 153854 118658
rect 153234 118338 153266 118574
rect 153502 118338 153586 118574
rect 153822 118338 153854 118574
rect 153234 82894 153854 118338
rect 153234 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 153854 82894
rect 153234 82574 153854 82658
rect 153234 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 153854 82574
rect 153234 46894 153854 82338
rect 153234 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 153854 46894
rect 153234 46574 153854 46658
rect 153234 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 153854 46574
rect 153234 10894 153854 46338
rect 153234 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 153854 10894
rect 153234 10574 153854 10658
rect 153234 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 153854 10574
rect 153234 -4186 153854 10338
rect 153234 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 153854 -4186
rect 153234 -4506 153854 -4422
rect 153234 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 153854 -4506
rect 153234 -5734 153854 -4742
rect 156954 194614 157574 198000
rect 156954 194378 156986 194614
rect 157222 194378 157306 194614
rect 157542 194378 157574 194614
rect 156954 194294 157574 194378
rect 156954 194058 156986 194294
rect 157222 194058 157306 194294
rect 157542 194058 157574 194294
rect 156954 158614 157574 194058
rect 156954 158378 156986 158614
rect 157222 158378 157306 158614
rect 157542 158378 157574 158614
rect 156954 158294 157574 158378
rect 156954 158058 156986 158294
rect 157222 158058 157306 158294
rect 157542 158058 157574 158294
rect 156954 122614 157574 158058
rect 156954 122378 156986 122614
rect 157222 122378 157306 122614
rect 157542 122378 157574 122614
rect 156954 122294 157574 122378
rect 156954 122058 156986 122294
rect 157222 122058 157306 122294
rect 157542 122058 157574 122294
rect 156954 86614 157574 122058
rect 156954 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 157574 86614
rect 156954 86294 157574 86378
rect 156954 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 157574 86294
rect 156954 50614 157574 86058
rect 156954 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 157574 50614
rect 156954 50294 157574 50378
rect 156954 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 157574 50294
rect 156954 14614 157574 50058
rect 156954 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 157574 14614
rect 156954 14294 157574 14378
rect 156954 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 157574 14294
rect 138954 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 139574 -7066
rect 138954 -7386 139574 -7302
rect 138954 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 139574 -7386
rect 138954 -7654 139574 -7622
rect 156954 -6106 157574 14058
rect 163794 165454 164414 198000
rect 163794 165218 163826 165454
rect 164062 165218 164146 165454
rect 164382 165218 164414 165454
rect 163794 165134 164414 165218
rect 163794 164898 163826 165134
rect 164062 164898 164146 165134
rect 164382 164898 164414 165134
rect 163794 129454 164414 164898
rect 163794 129218 163826 129454
rect 164062 129218 164146 129454
rect 164382 129218 164414 129454
rect 163794 129134 164414 129218
rect 163794 128898 163826 129134
rect 164062 128898 164146 129134
rect 164382 128898 164414 129134
rect 163794 93454 164414 128898
rect 163794 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 164414 93454
rect 163794 93134 164414 93218
rect 163794 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 164414 93134
rect 163794 57454 164414 92898
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -1306 164414 20898
rect 163794 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 164414 -1306
rect 163794 -1626 164414 -1542
rect 163794 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 164414 -1626
rect 163794 -1894 164414 -1862
rect 167514 169174 168134 198000
rect 167514 168938 167546 169174
rect 167782 168938 167866 169174
rect 168102 168938 168134 169174
rect 167514 168854 168134 168938
rect 167514 168618 167546 168854
rect 167782 168618 167866 168854
rect 168102 168618 168134 168854
rect 167514 133174 168134 168618
rect 167514 132938 167546 133174
rect 167782 132938 167866 133174
rect 168102 132938 168134 133174
rect 167514 132854 168134 132938
rect 167514 132618 167546 132854
rect 167782 132618 167866 132854
rect 168102 132618 168134 132854
rect 167514 97174 168134 132618
rect 167514 96938 167546 97174
rect 167782 96938 167866 97174
rect 168102 96938 168134 97174
rect 167514 96854 168134 96938
rect 167514 96618 167546 96854
rect 167782 96618 167866 96854
rect 168102 96618 168134 96854
rect 167514 61174 168134 96618
rect 167514 60938 167546 61174
rect 167782 60938 167866 61174
rect 168102 60938 168134 61174
rect 167514 60854 168134 60938
rect 167514 60618 167546 60854
rect 167782 60618 167866 60854
rect 168102 60618 168134 60854
rect 167514 25174 168134 60618
rect 167514 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 168134 25174
rect 167514 24854 168134 24938
rect 167514 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 168134 24854
rect 167514 -3226 168134 24618
rect 167514 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 168134 -3226
rect 167514 -3546 168134 -3462
rect 167514 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 168134 -3546
rect 167514 -3814 168134 -3782
rect 171234 172894 171854 198000
rect 173206 197845 173266 199550
rect 173390 198661 173450 199550
rect 173387 198660 173453 198661
rect 173387 198596 173388 198660
rect 173452 198596 173453 198660
rect 173387 198595 173453 198596
rect 186822 198117 186882 270539
rect 187003 234700 187069 234701
rect 187003 234636 187004 234700
rect 187068 234636 187069 234700
rect 187003 234635 187069 234636
rect 187006 198389 187066 234635
rect 187555 200700 187621 200701
rect 187555 200636 187556 200700
rect 187620 200636 187621 200700
rect 187555 200635 187621 200636
rect 187003 198388 187069 198389
rect 187003 198324 187004 198388
rect 187068 198324 187069 198388
rect 187003 198323 187069 198324
rect 187558 198253 187618 200635
rect 188294 199205 188354 285771
rect 189234 262894 189854 298338
rect 189234 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 189854 262894
rect 189234 262574 189854 262658
rect 189234 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 189854 262574
rect 189234 226894 189854 262338
rect 189234 226658 189266 226894
rect 189502 226658 189586 226894
rect 189822 226658 189854 226894
rect 189234 226574 189854 226658
rect 189234 226338 189266 226574
rect 189502 226338 189586 226574
rect 189822 226338 189854 226574
rect 188475 222868 188541 222869
rect 188475 222804 188476 222868
rect 188540 222804 188541 222868
rect 188475 222803 188541 222804
rect 188291 199204 188357 199205
rect 188291 199140 188292 199204
rect 188356 199140 188357 199204
rect 188291 199139 188357 199140
rect 187555 198252 187621 198253
rect 187555 198188 187556 198252
rect 187620 198188 187621 198252
rect 187555 198187 187621 198188
rect 186819 198116 186885 198117
rect 186819 198052 186820 198116
rect 186884 198052 186885 198116
rect 186819 198051 186885 198052
rect 173203 197844 173269 197845
rect 173203 197780 173204 197844
rect 173268 197780 173269 197844
rect 173203 197779 173269 197780
rect 171234 172658 171266 172894
rect 171502 172658 171586 172894
rect 171822 172658 171854 172894
rect 171234 172574 171854 172658
rect 171234 172338 171266 172574
rect 171502 172338 171586 172574
rect 171822 172338 171854 172574
rect 171234 136894 171854 172338
rect 171234 136658 171266 136894
rect 171502 136658 171586 136894
rect 171822 136658 171854 136894
rect 171234 136574 171854 136658
rect 171234 136338 171266 136574
rect 171502 136338 171586 136574
rect 171822 136338 171854 136574
rect 171234 100894 171854 136338
rect 171234 100658 171266 100894
rect 171502 100658 171586 100894
rect 171822 100658 171854 100894
rect 171234 100574 171854 100658
rect 171234 100338 171266 100574
rect 171502 100338 171586 100574
rect 171822 100338 171854 100574
rect 171234 64894 171854 100338
rect 171234 64658 171266 64894
rect 171502 64658 171586 64894
rect 171822 64658 171854 64894
rect 171234 64574 171854 64658
rect 171234 64338 171266 64574
rect 171502 64338 171586 64574
rect 171822 64338 171854 64574
rect 171234 28894 171854 64338
rect 171234 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 171854 28894
rect 171234 28574 171854 28658
rect 171234 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 171854 28574
rect 171234 -5146 171854 28338
rect 171234 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 171854 -5146
rect 171234 -5466 171854 -5382
rect 171234 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 171854 -5466
rect 171234 -5734 171854 -5702
rect 174954 176614 175574 198000
rect 174954 176378 174986 176614
rect 175222 176378 175306 176614
rect 175542 176378 175574 176614
rect 174954 176294 175574 176378
rect 174954 176058 174986 176294
rect 175222 176058 175306 176294
rect 175542 176058 175574 176294
rect 174954 140614 175574 176058
rect 174954 140378 174986 140614
rect 175222 140378 175306 140614
rect 175542 140378 175574 140614
rect 174954 140294 175574 140378
rect 174954 140058 174986 140294
rect 175222 140058 175306 140294
rect 175542 140058 175574 140294
rect 174954 104614 175574 140058
rect 174954 104378 174986 104614
rect 175222 104378 175306 104614
rect 175542 104378 175574 104614
rect 174954 104294 175574 104378
rect 174954 104058 174986 104294
rect 175222 104058 175306 104294
rect 175542 104058 175574 104294
rect 174954 68614 175574 104058
rect 174954 68378 174986 68614
rect 175222 68378 175306 68614
rect 175542 68378 175574 68614
rect 174954 68294 175574 68378
rect 174954 68058 174986 68294
rect 175222 68058 175306 68294
rect 175542 68058 175574 68294
rect 174954 32614 175574 68058
rect 174954 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 175574 32614
rect 174954 32294 175574 32378
rect 174954 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 175574 32294
rect 156954 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 157574 -6106
rect 156954 -6426 157574 -6342
rect 156954 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 157574 -6426
rect 156954 -7654 157574 -6662
rect 174954 -7066 175574 32058
rect 181794 183454 182414 198000
rect 181794 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 182414 183454
rect 181794 183134 182414 183218
rect 181794 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 182414 183134
rect 181794 147454 182414 182898
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 111454 182414 146898
rect 181794 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 182414 111454
rect 181794 111134 182414 111218
rect 181794 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 182414 111134
rect 181794 75454 182414 110898
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 181794 39454 182414 74898
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -1894 182414 -902
rect 185514 187174 186134 198000
rect 188478 197981 188538 222803
rect 188475 197980 188541 197981
rect 188475 197916 188476 197980
rect 188540 197916 188541 197980
rect 188475 197915 188541 197916
rect 185514 186938 185546 187174
rect 185782 186938 185866 187174
rect 186102 186938 186134 187174
rect 185514 186854 186134 186938
rect 185514 186618 185546 186854
rect 185782 186618 185866 186854
rect 186102 186618 186134 186854
rect 185514 151174 186134 186618
rect 185514 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 186134 151174
rect 185514 150854 186134 150938
rect 185514 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 186134 150854
rect 185514 115174 186134 150618
rect 185514 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 186134 115174
rect 185514 114854 186134 114938
rect 185514 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 186134 114854
rect 185514 79174 186134 114618
rect 185514 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 186134 79174
rect 185514 78854 186134 78938
rect 185514 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 186134 78854
rect 185514 43174 186134 78618
rect 185514 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 186134 43174
rect 185514 42854 186134 42938
rect 185514 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 186134 42854
rect 185514 7174 186134 42618
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 185514 -2266 186134 6618
rect 185514 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 186134 -2266
rect 185514 -2586 186134 -2502
rect 185514 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 186134 -2586
rect 185514 -3814 186134 -2822
rect 189234 190894 189854 226338
rect 189234 190658 189266 190894
rect 189502 190658 189586 190894
rect 189822 190658 189854 190894
rect 189234 190574 189854 190658
rect 189234 190338 189266 190574
rect 189502 190338 189586 190574
rect 189822 190338 189854 190574
rect 189234 154894 189854 190338
rect 189234 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 189854 154894
rect 189234 154574 189854 154658
rect 189234 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 189854 154574
rect 189234 118894 189854 154338
rect 189234 118658 189266 118894
rect 189502 118658 189586 118894
rect 189822 118658 189854 118894
rect 189234 118574 189854 118658
rect 189234 118338 189266 118574
rect 189502 118338 189586 118574
rect 189822 118338 189854 118574
rect 189234 82894 189854 118338
rect 189234 82658 189266 82894
rect 189502 82658 189586 82894
rect 189822 82658 189854 82894
rect 189234 82574 189854 82658
rect 189234 82338 189266 82574
rect 189502 82338 189586 82574
rect 189822 82338 189854 82574
rect 189234 46894 189854 82338
rect 189234 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 189854 46894
rect 189234 46574 189854 46658
rect 189234 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 189854 46574
rect 189234 10894 189854 46338
rect 189234 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 189854 10894
rect 189234 10574 189854 10658
rect 189234 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 189854 10574
rect 189234 -4186 189854 10338
rect 189234 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 189854 -4186
rect 189234 -4506 189854 -4422
rect 189234 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 189854 -4506
rect 189234 -5734 189854 -4742
rect 192954 698614 193574 710042
rect 210954 711558 211574 711590
rect 210954 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 211574 711558
rect 210954 711238 211574 711322
rect 210954 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 211574 711238
rect 207234 709638 207854 709670
rect 207234 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 207854 709638
rect 207234 709318 207854 709402
rect 207234 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 207854 709318
rect 203514 707718 204134 707750
rect 203514 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 204134 707718
rect 203514 707398 204134 707482
rect 203514 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 204134 707398
rect 192954 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 193574 698614
rect 192954 698294 193574 698378
rect 192954 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 193574 698294
rect 192954 662614 193574 698058
rect 192954 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 193574 662614
rect 192954 662294 193574 662378
rect 192954 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 193574 662294
rect 192954 626614 193574 662058
rect 192954 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 193574 626614
rect 192954 626294 193574 626378
rect 192954 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 193574 626294
rect 192954 590614 193574 626058
rect 192954 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 193574 590614
rect 192954 590294 193574 590378
rect 192954 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 193574 590294
rect 192954 554614 193574 590058
rect 192954 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 193574 554614
rect 192954 554294 193574 554378
rect 192954 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 193574 554294
rect 192954 518614 193574 554058
rect 192954 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 193574 518614
rect 192954 518294 193574 518378
rect 192954 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 193574 518294
rect 192954 482614 193574 518058
rect 192954 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 193574 482614
rect 192954 482294 193574 482378
rect 192954 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 193574 482294
rect 192954 446614 193574 482058
rect 192954 446378 192986 446614
rect 193222 446378 193306 446614
rect 193542 446378 193574 446614
rect 192954 446294 193574 446378
rect 192954 446058 192986 446294
rect 193222 446058 193306 446294
rect 193542 446058 193574 446294
rect 192954 410614 193574 446058
rect 192954 410378 192986 410614
rect 193222 410378 193306 410614
rect 193542 410378 193574 410614
rect 192954 410294 193574 410378
rect 192954 410058 192986 410294
rect 193222 410058 193306 410294
rect 193542 410058 193574 410294
rect 192954 374614 193574 410058
rect 192954 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 193574 374614
rect 192954 374294 193574 374378
rect 192954 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 193574 374294
rect 192954 338614 193574 374058
rect 192954 338378 192986 338614
rect 193222 338378 193306 338614
rect 193542 338378 193574 338614
rect 192954 338294 193574 338378
rect 192954 338058 192986 338294
rect 193222 338058 193306 338294
rect 193542 338058 193574 338294
rect 192954 302614 193574 338058
rect 192954 302378 192986 302614
rect 193222 302378 193306 302614
rect 193542 302378 193574 302614
rect 192954 302294 193574 302378
rect 192954 302058 192986 302294
rect 193222 302058 193306 302294
rect 193542 302058 193574 302294
rect 192954 266614 193574 302058
rect 192954 266378 192986 266614
rect 193222 266378 193306 266614
rect 193542 266378 193574 266614
rect 192954 266294 193574 266378
rect 192954 266058 192986 266294
rect 193222 266058 193306 266294
rect 193542 266058 193574 266294
rect 192954 230614 193574 266058
rect 192954 230378 192986 230614
rect 193222 230378 193306 230614
rect 193542 230378 193574 230614
rect 192954 230294 193574 230378
rect 192954 230058 192986 230294
rect 193222 230058 193306 230294
rect 193542 230058 193574 230294
rect 192954 194614 193574 230058
rect 192954 194378 192986 194614
rect 193222 194378 193306 194614
rect 193542 194378 193574 194614
rect 192954 194294 193574 194378
rect 192954 194058 192986 194294
rect 193222 194058 193306 194294
rect 193542 194058 193574 194294
rect 192954 158614 193574 194058
rect 192954 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 193574 158614
rect 192954 158294 193574 158378
rect 192954 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 193574 158294
rect 192954 122614 193574 158058
rect 192954 122378 192986 122614
rect 193222 122378 193306 122614
rect 193542 122378 193574 122614
rect 192954 122294 193574 122378
rect 192954 122058 192986 122294
rect 193222 122058 193306 122294
rect 193542 122058 193574 122294
rect 192954 86614 193574 122058
rect 192954 86378 192986 86614
rect 193222 86378 193306 86614
rect 193542 86378 193574 86614
rect 192954 86294 193574 86378
rect 192954 86058 192986 86294
rect 193222 86058 193306 86294
rect 193542 86058 193574 86294
rect 192954 50614 193574 86058
rect 192954 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 193574 50614
rect 192954 50294 193574 50378
rect 192954 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 193574 50294
rect 192954 14614 193574 50058
rect 192954 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 193574 14614
rect 192954 14294 193574 14378
rect 192954 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 193574 14294
rect 174954 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 175574 -7066
rect 174954 -7386 175574 -7302
rect 174954 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 175574 -7386
rect 174954 -7654 175574 -7622
rect 192954 -6106 193574 14058
rect 199794 705798 200414 705830
rect 199794 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 200414 705798
rect 199794 705478 200414 705562
rect 199794 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 200414 705478
rect 199794 669454 200414 705242
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 561454 200414 596898
rect 199794 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 200414 561454
rect 199794 561134 200414 561218
rect 199794 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 200414 561134
rect 199794 525454 200414 560898
rect 199794 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 200414 525454
rect 199794 525134 200414 525218
rect 199794 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 200414 525134
rect 199794 489454 200414 524898
rect 199794 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 200414 489454
rect 199794 489134 200414 489218
rect 199794 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 200414 489134
rect 199794 453454 200414 488898
rect 199794 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 200414 453454
rect 199794 453134 200414 453218
rect 199794 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 200414 453134
rect 199794 417454 200414 452898
rect 199794 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 200414 417454
rect 199794 417134 200414 417218
rect 199794 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 200414 417134
rect 199794 381454 200414 416898
rect 199794 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 200414 381454
rect 199794 381134 200414 381218
rect 199794 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 200414 381134
rect 199794 345454 200414 380898
rect 199794 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 200414 345454
rect 199794 345134 200414 345218
rect 199794 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 200414 345134
rect 199794 309454 200414 344898
rect 199794 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 200414 309454
rect 199794 309134 200414 309218
rect 199794 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 200414 309134
rect 199794 273454 200414 308898
rect 199794 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 200414 273454
rect 199794 273134 200414 273218
rect 199794 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 200414 273134
rect 199794 237454 200414 272898
rect 199794 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 200414 237454
rect 199794 237134 200414 237218
rect 199794 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 200414 237134
rect 199794 201454 200414 236898
rect 199794 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 200414 201454
rect 199794 201134 200414 201218
rect 199794 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 200414 201134
rect 199794 165454 200414 200898
rect 199794 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 200414 165454
rect 199794 165134 200414 165218
rect 199794 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 200414 165134
rect 199794 129454 200414 164898
rect 199794 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 200414 129454
rect 199794 129134 200414 129218
rect 199794 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 200414 129134
rect 199794 93454 200414 128898
rect 199794 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 200414 93454
rect 199794 93134 200414 93218
rect 199794 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 200414 93134
rect 199794 57454 200414 92898
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -1306 200414 20898
rect 199794 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 200414 -1306
rect 199794 -1626 200414 -1542
rect 199794 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 200414 -1626
rect 199794 -1894 200414 -1862
rect 203514 673174 204134 707162
rect 203514 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 204134 673174
rect 203514 672854 204134 672938
rect 203514 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 204134 672854
rect 203514 637174 204134 672618
rect 203514 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 204134 637174
rect 203514 636854 204134 636938
rect 203514 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 204134 636854
rect 203514 601174 204134 636618
rect 203514 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 204134 601174
rect 203514 600854 204134 600938
rect 203514 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 204134 600854
rect 203514 565174 204134 600618
rect 203514 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 204134 565174
rect 203514 564854 204134 564938
rect 203514 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 204134 564854
rect 203514 529174 204134 564618
rect 203514 528938 203546 529174
rect 203782 528938 203866 529174
rect 204102 528938 204134 529174
rect 203514 528854 204134 528938
rect 203514 528618 203546 528854
rect 203782 528618 203866 528854
rect 204102 528618 204134 528854
rect 203514 493174 204134 528618
rect 203514 492938 203546 493174
rect 203782 492938 203866 493174
rect 204102 492938 204134 493174
rect 203514 492854 204134 492938
rect 203514 492618 203546 492854
rect 203782 492618 203866 492854
rect 204102 492618 204134 492854
rect 203514 457174 204134 492618
rect 203514 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 204134 457174
rect 203514 456854 204134 456938
rect 203514 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 204134 456854
rect 203514 421174 204134 456618
rect 203514 420938 203546 421174
rect 203782 420938 203866 421174
rect 204102 420938 204134 421174
rect 203514 420854 204134 420938
rect 203514 420618 203546 420854
rect 203782 420618 203866 420854
rect 204102 420618 204134 420854
rect 203514 385174 204134 420618
rect 203514 384938 203546 385174
rect 203782 384938 203866 385174
rect 204102 384938 204134 385174
rect 203514 384854 204134 384938
rect 203514 384618 203546 384854
rect 203782 384618 203866 384854
rect 204102 384618 204134 384854
rect 203514 349174 204134 384618
rect 203514 348938 203546 349174
rect 203782 348938 203866 349174
rect 204102 348938 204134 349174
rect 203514 348854 204134 348938
rect 203514 348618 203546 348854
rect 203782 348618 203866 348854
rect 204102 348618 204134 348854
rect 203514 313174 204134 348618
rect 203514 312938 203546 313174
rect 203782 312938 203866 313174
rect 204102 312938 204134 313174
rect 203514 312854 204134 312938
rect 203514 312618 203546 312854
rect 203782 312618 203866 312854
rect 204102 312618 204134 312854
rect 203514 277174 204134 312618
rect 203514 276938 203546 277174
rect 203782 276938 203866 277174
rect 204102 276938 204134 277174
rect 203514 276854 204134 276938
rect 203514 276618 203546 276854
rect 203782 276618 203866 276854
rect 204102 276618 204134 276854
rect 203514 241174 204134 276618
rect 203514 240938 203546 241174
rect 203782 240938 203866 241174
rect 204102 240938 204134 241174
rect 203514 240854 204134 240938
rect 203514 240618 203546 240854
rect 203782 240618 203866 240854
rect 204102 240618 204134 240854
rect 203514 205174 204134 240618
rect 203514 204938 203546 205174
rect 203782 204938 203866 205174
rect 204102 204938 204134 205174
rect 203514 204854 204134 204938
rect 203514 204618 203546 204854
rect 203782 204618 203866 204854
rect 204102 204618 204134 204854
rect 203514 169174 204134 204618
rect 203514 168938 203546 169174
rect 203782 168938 203866 169174
rect 204102 168938 204134 169174
rect 203514 168854 204134 168938
rect 203514 168618 203546 168854
rect 203782 168618 203866 168854
rect 204102 168618 204134 168854
rect 203514 133174 204134 168618
rect 203514 132938 203546 133174
rect 203782 132938 203866 133174
rect 204102 132938 204134 133174
rect 203514 132854 204134 132938
rect 203514 132618 203546 132854
rect 203782 132618 203866 132854
rect 204102 132618 204134 132854
rect 203514 97174 204134 132618
rect 203514 96938 203546 97174
rect 203782 96938 203866 97174
rect 204102 96938 204134 97174
rect 203514 96854 204134 96938
rect 203514 96618 203546 96854
rect 203782 96618 203866 96854
rect 204102 96618 204134 96854
rect 203514 61174 204134 96618
rect 203514 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 204134 61174
rect 203514 60854 204134 60938
rect 203514 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 204134 60854
rect 203514 25174 204134 60618
rect 203514 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 204134 25174
rect 203514 24854 204134 24938
rect 203514 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 204134 24854
rect 203514 -3226 204134 24618
rect 203514 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 204134 -3226
rect 203514 -3546 204134 -3462
rect 203514 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 204134 -3546
rect 203514 -3814 204134 -3782
rect 207234 676894 207854 709082
rect 207234 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 207854 676894
rect 207234 676574 207854 676658
rect 207234 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 207854 676574
rect 207234 640894 207854 676338
rect 207234 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 207854 640894
rect 207234 640574 207854 640658
rect 207234 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 207854 640574
rect 207234 604894 207854 640338
rect 207234 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 207854 604894
rect 207234 604574 207854 604658
rect 207234 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 207854 604574
rect 207234 568894 207854 604338
rect 207234 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 207854 568894
rect 207234 568574 207854 568658
rect 207234 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 207854 568574
rect 207234 532894 207854 568338
rect 207234 532658 207266 532894
rect 207502 532658 207586 532894
rect 207822 532658 207854 532894
rect 207234 532574 207854 532658
rect 207234 532338 207266 532574
rect 207502 532338 207586 532574
rect 207822 532338 207854 532574
rect 207234 496894 207854 532338
rect 207234 496658 207266 496894
rect 207502 496658 207586 496894
rect 207822 496658 207854 496894
rect 207234 496574 207854 496658
rect 207234 496338 207266 496574
rect 207502 496338 207586 496574
rect 207822 496338 207854 496574
rect 207234 460894 207854 496338
rect 207234 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 207854 460894
rect 207234 460574 207854 460658
rect 207234 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 207854 460574
rect 207234 424894 207854 460338
rect 207234 424658 207266 424894
rect 207502 424658 207586 424894
rect 207822 424658 207854 424894
rect 207234 424574 207854 424658
rect 207234 424338 207266 424574
rect 207502 424338 207586 424574
rect 207822 424338 207854 424574
rect 207234 388894 207854 424338
rect 207234 388658 207266 388894
rect 207502 388658 207586 388894
rect 207822 388658 207854 388894
rect 207234 388574 207854 388658
rect 207234 388338 207266 388574
rect 207502 388338 207586 388574
rect 207822 388338 207854 388574
rect 207234 352894 207854 388338
rect 207234 352658 207266 352894
rect 207502 352658 207586 352894
rect 207822 352658 207854 352894
rect 207234 352574 207854 352658
rect 207234 352338 207266 352574
rect 207502 352338 207586 352574
rect 207822 352338 207854 352574
rect 207234 316894 207854 352338
rect 207234 316658 207266 316894
rect 207502 316658 207586 316894
rect 207822 316658 207854 316894
rect 207234 316574 207854 316658
rect 207234 316338 207266 316574
rect 207502 316338 207586 316574
rect 207822 316338 207854 316574
rect 207234 280894 207854 316338
rect 207234 280658 207266 280894
rect 207502 280658 207586 280894
rect 207822 280658 207854 280894
rect 207234 280574 207854 280658
rect 207234 280338 207266 280574
rect 207502 280338 207586 280574
rect 207822 280338 207854 280574
rect 207234 244894 207854 280338
rect 207234 244658 207266 244894
rect 207502 244658 207586 244894
rect 207822 244658 207854 244894
rect 207234 244574 207854 244658
rect 207234 244338 207266 244574
rect 207502 244338 207586 244574
rect 207822 244338 207854 244574
rect 207234 208894 207854 244338
rect 207234 208658 207266 208894
rect 207502 208658 207586 208894
rect 207822 208658 207854 208894
rect 207234 208574 207854 208658
rect 207234 208338 207266 208574
rect 207502 208338 207586 208574
rect 207822 208338 207854 208574
rect 207234 172894 207854 208338
rect 207234 172658 207266 172894
rect 207502 172658 207586 172894
rect 207822 172658 207854 172894
rect 207234 172574 207854 172658
rect 207234 172338 207266 172574
rect 207502 172338 207586 172574
rect 207822 172338 207854 172574
rect 207234 136894 207854 172338
rect 207234 136658 207266 136894
rect 207502 136658 207586 136894
rect 207822 136658 207854 136894
rect 207234 136574 207854 136658
rect 207234 136338 207266 136574
rect 207502 136338 207586 136574
rect 207822 136338 207854 136574
rect 207234 100894 207854 136338
rect 207234 100658 207266 100894
rect 207502 100658 207586 100894
rect 207822 100658 207854 100894
rect 207234 100574 207854 100658
rect 207234 100338 207266 100574
rect 207502 100338 207586 100574
rect 207822 100338 207854 100574
rect 207234 64894 207854 100338
rect 207234 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 207854 64894
rect 207234 64574 207854 64658
rect 207234 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 207854 64574
rect 207234 28894 207854 64338
rect 207234 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 207854 28894
rect 207234 28574 207854 28658
rect 207234 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 207854 28574
rect 207234 -5146 207854 28338
rect 207234 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 207854 -5146
rect 207234 -5466 207854 -5382
rect 207234 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 207854 -5466
rect 207234 -5734 207854 -5702
rect 210954 680614 211574 711002
rect 228954 710598 229574 711590
rect 228954 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 229574 710598
rect 228954 710278 229574 710362
rect 228954 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 229574 710278
rect 225234 708678 225854 709670
rect 225234 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 225854 708678
rect 225234 708358 225854 708442
rect 225234 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 225854 708358
rect 221514 706758 222134 707750
rect 221514 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 222134 706758
rect 221514 706438 222134 706522
rect 221514 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 222134 706438
rect 210954 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 211574 680614
rect 210954 680294 211574 680378
rect 210954 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 211574 680294
rect 210954 644614 211574 680058
rect 210954 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 211574 644614
rect 210954 644294 211574 644378
rect 210954 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 211574 644294
rect 210954 608614 211574 644058
rect 210954 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 211574 608614
rect 210954 608294 211574 608378
rect 210954 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 211574 608294
rect 210954 572614 211574 608058
rect 210954 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 211574 572614
rect 210954 572294 211574 572378
rect 210954 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 211574 572294
rect 210954 536614 211574 572058
rect 210954 536378 210986 536614
rect 211222 536378 211306 536614
rect 211542 536378 211574 536614
rect 210954 536294 211574 536378
rect 210954 536058 210986 536294
rect 211222 536058 211306 536294
rect 211542 536058 211574 536294
rect 210954 500614 211574 536058
rect 210954 500378 210986 500614
rect 211222 500378 211306 500614
rect 211542 500378 211574 500614
rect 210954 500294 211574 500378
rect 210954 500058 210986 500294
rect 211222 500058 211306 500294
rect 211542 500058 211574 500294
rect 210954 464614 211574 500058
rect 210954 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 211574 464614
rect 210954 464294 211574 464378
rect 210954 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 211574 464294
rect 210954 428614 211574 464058
rect 210954 428378 210986 428614
rect 211222 428378 211306 428614
rect 211542 428378 211574 428614
rect 210954 428294 211574 428378
rect 210954 428058 210986 428294
rect 211222 428058 211306 428294
rect 211542 428058 211574 428294
rect 210954 392614 211574 428058
rect 210954 392378 210986 392614
rect 211222 392378 211306 392614
rect 211542 392378 211574 392614
rect 210954 392294 211574 392378
rect 210954 392058 210986 392294
rect 211222 392058 211306 392294
rect 211542 392058 211574 392294
rect 210954 356614 211574 392058
rect 210954 356378 210986 356614
rect 211222 356378 211306 356614
rect 211542 356378 211574 356614
rect 210954 356294 211574 356378
rect 210954 356058 210986 356294
rect 211222 356058 211306 356294
rect 211542 356058 211574 356294
rect 210954 320614 211574 356058
rect 210954 320378 210986 320614
rect 211222 320378 211306 320614
rect 211542 320378 211574 320614
rect 210954 320294 211574 320378
rect 210954 320058 210986 320294
rect 211222 320058 211306 320294
rect 211542 320058 211574 320294
rect 210954 284614 211574 320058
rect 210954 284378 210986 284614
rect 211222 284378 211306 284614
rect 211542 284378 211574 284614
rect 210954 284294 211574 284378
rect 210954 284058 210986 284294
rect 211222 284058 211306 284294
rect 211542 284058 211574 284294
rect 210954 248614 211574 284058
rect 210954 248378 210986 248614
rect 211222 248378 211306 248614
rect 211542 248378 211574 248614
rect 210954 248294 211574 248378
rect 210954 248058 210986 248294
rect 211222 248058 211306 248294
rect 211542 248058 211574 248294
rect 210954 212614 211574 248058
rect 210954 212378 210986 212614
rect 211222 212378 211306 212614
rect 211542 212378 211574 212614
rect 210954 212294 211574 212378
rect 210954 212058 210986 212294
rect 211222 212058 211306 212294
rect 211542 212058 211574 212294
rect 210954 176614 211574 212058
rect 210954 176378 210986 176614
rect 211222 176378 211306 176614
rect 211542 176378 211574 176614
rect 210954 176294 211574 176378
rect 210954 176058 210986 176294
rect 211222 176058 211306 176294
rect 211542 176058 211574 176294
rect 210954 140614 211574 176058
rect 210954 140378 210986 140614
rect 211222 140378 211306 140614
rect 211542 140378 211574 140614
rect 210954 140294 211574 140378
rect 210954 140058 210986 140294
rect 211222 140058 211306 140294
rect 211542 140058 211574 140294
rect 210954 104614 211574 140058
rect 210954 104378 210986 104614
rect 211222 104378 211306 104614
rect 211542 104378 211574 104614
rect 210954 104294 211574 104378
rect 210954 104058 210986 104294
rect 211222 104058 211306 104294
rect 211542 104058 211574 104294
rect 210954 68614 211574 104058
rect 210954 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 211574 68614
rect 210954 68294 211574 68378
rect 210954 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 211574 68294
rect 210954 32614 211574 68058
rect 210954 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 211574 32614
rect 210954 32294 211574 32378
rect 210954 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 211574 32294
rect 192954 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 193574 -6106
rect 192954 -6426 193574 -6342
rect 192954 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 193574 -6426
rect 192954 -7654 193574 -6662
rect 210954 -7066 211574 32058
rect 217794 704838 218414 705830
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 543454 218414 578898
rect 217794 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 218414 543454
rect 217794 543134 218414 543218
rect 217794 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 218414 543134
rect 217794 507454 218414 542898
rect 217794 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 218414 507454
rect 217794 507134 218414 507218
rect 217794 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 218414 507134
rect 217794 471454 218414 506898
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 217794 435454 218414 470898
rect 217794 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 218414 435454
rect 217794 435134 218414 435218
rect 217794 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 218414 435134
rect 217794 399454 218414 434898
rect 217794 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 218414 399454
rect 217794 399134 218414 399218
rect 217794 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 218414 399134
rect 217794 363454 218414 398898
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 217794 327454 218414 362898
rect 217794 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 218414 327454
rect 217794 327134 218414 327218
rect 217794 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 218414 327134
rect 217794 291454 218414 326898
rect 217794 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 218414 291454
rect 217794 291134 218414 291218
rect 217794 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 218414 291134
rect 217794 255454 218414 290898
rect 217794 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 218414 255454
rect 217794 255134 218414 255218
rect 217794 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 218414 255134
rect 217794 219454 218414 254898
rect 217794 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 218414 219454
rect 217794 219134 218414 219218
rect 217794 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 218414 219134
rect 217794 183454 218414 218898
rect 217794 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 218414 183454
rect 217794 183134 218414 183218
rect 217794 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 218414 183134
rect 217794 147454 218414 182898
rect 217794 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 218414 147454
rect 217794 147134 218414 147218
rect 217794 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 218414 147134
rect 217794 111454 218414 146898
rect 217794 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 218414 111454
rect 217794 111134 218414 111218
rect 217794 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 218414 111134
rect 217794 75454 218414 110898
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 217794 39454 218414 74898
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -1894 218414 -902
rect 221514 691174 222134 706202
rect 221514 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 222134 691174
rect 221514 690854 222134 690938
rect 221514 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 222134 690854
rect 221514 655174 222134 690618
rect 221514 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 222134 655174
rect 221514 654854 222134 654938
rect 221514 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 222134 654854
rect 221514 619174 222134 654618
rect 221514 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 222134 619174
rect 221514 618854 222134 618938
rect 221514 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 222134 618854
rect 221514 583174 222134 618618
rect 221514 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 222134 583174
rect 221514 582854 222134 582938
rect 221514 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 222134 582854
rect 221514 547174 222134 582618
rect 221514 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 222134 547174
rect 221514 546854 222134 546938
rect 221514 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 222134 546854
rect 221514 511174 222134 546618
rect 221514 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 222134 511174
rect 221514 510854 222134 510938
rect 221514 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 222134 510854
rect 221514 475174 222134 510618
rect 221514 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 222134 475174
rect 221514 474854 222134 474938
rect 221514 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 222134 474854
rect 221514 439174 222134 474618
rect 221514 438938 221546 439174
rect 221782 438938 221866 439174
rect 222102 438938 222134 439174
rect 221514 438854 222134 438938
rect 221514 438618 221546 438854
rect 221782 438618 221866 438854
rect 222102 438618 222134 438854
rect 221514 403174 222134 438618
rect 221514 402938 221546 403174
rect 221782 402938 221866 403174
rect 222102 402938 222134 403174
rect 221514 402854 222134 402938
rect 221514 402618 221546 402854
rect 221782 402618 221866 402854
rect 222102 402618 222134 402854
rect 221514 367174 222134 402618
rect 221514 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 222134 367174
rect 221514 366854 222134 366938
rect 221514 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 222134 366854
rect 221514 331174 222134 366618
rect 221514 330938 221546 331174
rect 221782 330938 221866 331174
rect 222102 330938 222134 331174
rect 221514 330854 222134 330938
rect 221514 330618 221546 330854
rect 221782 330618 221866 330854
rect 222102 330618 222134 330854
rect 221514 295174 222134 330618
rect 221514 294938 221546 295174
rect 221782 294938 221866 295174
rect 222102 294938 222134 295174
rect 221514 294854 222134 294938
rect 221514 294618 221546 294854
rect 221782 294618 221866 294854
rect 222102 294618 222134 294854
rect 221514 259174 222134 294618
rect 221514 258938 221546 259174
rect 221782 258938 221866 259174
rect 222102 258938 222134 259174
rect 221514 258854 222134 258938
rect 221514 258618 221546 258854
rect 221782 258618 221866 258854
rect 222102 258618 222134 258854
rect 221514 223174 222134 258618
rect 221514 222938 221546 223174
rect 221782 222938 221866 223174
rect 222102 222938 222134 223174
rect 221514 222854 222134 222938
rect 221514 222618 221546 222854
rect 221782 222618 221866 222854
rect 222102 222618 222134 222854
rect 221514 187174 222134 222618
rect 221514 186938 221546 187174
rect 221782 186938 221866 187174
rect 222102 186938 222134 187174
rect 221514 186854 222134 186938
rect 221514 186618 221546 186854
rect 221782 186618 221866 186854
rect 222102 186618 222134 186854
rect 221514 151174 222134 186618
rect 221514 150938 221546 151174
rect 221782 150938 221866 151174
rect 222102 150938 222134 151174
rect 221514 150854 222134 150938
rect 221514 150618 221546 150854
rect 221782 150618 221866 150854
rect 222102 150618 222134 150854
rect 221514 115174 222134 150618
rect 221514 114938 221546 115174
rect 221782 114938 221866 115174
rect 222102 114938 222134 115174
rect 221514 114854 222134 114938
rect 221514 114618 221546 114854
rect 221782 114618 221866 114854
rect 222102 114618 222134 114854
rect 221514 79174 222134 114618
rect 221514 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 222134 79174
rect 221514 78854 222134 78938
rect 221514 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 222134 78854
rect 221514 43174 222134 78618
rect 221514 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 222134 43174
rect 221514 42854 222134 42938
rect 221514 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 222134 42854
rect 221514 7174 222134 42618
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -2266 222134 6618
rect 221514 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 222134 -2266
rect 221514 -2586 222134 -2502
rect 221514 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 222134 -2586
rect 221514 -3814 222134 -2822
rect 225234 694894 225854 708122
rect 225234 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 225854 694894
rect 225234 694574 225854 694658
rect 225234 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 225854 694574
rect 225234 658894 225854 694338
rect 225234 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 225854 658894
rect 225234 658574 225854 658658
rect 225234 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 225854 658574
rect 225234 622894 225854 658338
rect 225234 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 225854 622894
rect 225234 622574 225854 622658
rect 225234 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 225854 622574
rect 225234 586894 225854 622338
rect 225234 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 225854 586894
rect 225234 586574 225854 586658
rect 225234 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 225854 586574
rect 225234 550894 225854 586338
rect 225234 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 225854 550894
rect 225234 550574 225854 550658
rect 225234 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 225854 550574
rect 225234 514894 225854 550338
rect 225234 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 225854 514894
rect 225234 514574 225854 514658
rect 225234 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 225854 514574
rect 225234 478894 225854 514338
rect 225234 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 225854 478894
rect 225234 478574 225854 478658
rect 225234 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 225854 478574
rect 225234 442894 225854 478338
rect 225234 442658 225266 442894
rect 225502 442658 225586 442894
rect 225822 442658 225854 442894
rect 225234 442574 225854 442658
rect 225234 442338 225266 442574
rect 225502 442338 225586 442574
rect 225822 442338 225854 442574
rect 225234 406894 225854 442338
rect 225234 406658 225266 406894
rect 225502 406658 225586 406894
rect 225822 406658 225854 406894
rect 225234 406574 225854 406658
rect 225234 406338 225266 406574
rect 225502 406338 225586 406574
rect 225822 406338 225854 406574
rect 225234 370894 225854 406338
rect 225234 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 225854 370894
rect 225234 370574 225854 370658
rect 225234 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 225854 370574
rect 225234 334894 225854 370338
rect 225234 334658 225266 334894
rect 225502 334658 225586 334894
rect 225822 334658 225854 334894
rect 225234 334574 225854 334658
rect 225234 334338 225266 334574
rect 225502 334338 225586 334574
rect 225822 334338 225854 334574
rect 225234 298894 225854 334338
rect 225234 298658 225266 298894
rect 225502 298658 225586 298894
rect 225822 298658 225854 298894
rect 225234 298574 225854 298658
rect 225234 298338 225266 298574
rect 225502 298338 225586 298574
rect 225822 298338 225854 298574
rect 225234 262894 225854 298338
rect 225234 262658 225266 262894
rect 225502 262658 225586 262894
rect 225822 262658 225854 262894
rect 225234 262574 225854 262658
rect 225234 262338 225266 262574
rect 225502 262338 225586 262574
rect 225822 262338 225854 262574
rect 225234 226894 225854 262338
rect 225234 226658 225266 226894
rect 225502 226658 225586 226894
rect 225822 226658 225854 226894
rect 225234 226574 225854 226658
rect 225234 226338 225266 226574
rect 225502 226338 225586 226574
rect 225822 226338 225854 226574
rect 225234 190894 225854 226338
rect 225234 190658 225266 190894
rect 225502 190658 225586 190894
rect 225822 190658 225854 190894
rect 225234 190574 225854 190658
rect 225234 190338 225266 190574
rect 225502 190338 225586 190574
rect 225822 190338 225854 190574
rect 225234 154894 225854 190338
rect 225234 154658 225266 154894
rect 225502 154658 225586 154894
rect 225822 154658 225854 154894
rect 225234 154574 225854 154658
rect 225234 154338 225266 154574
rect 225502 154338 225586 154574
rect 225822 154338 225854 154574
rect 225234 118894 225854 154338
rect 225234 118658 225266 118894
rect 225502 118658 225586 118894
rect 225822 118658 225854 118894
rect 225234 118574 225854 118658
rect 225234 118338 225266 118574
rect 225502 118338 225586 118574
rect 225822 118338 225854 118574
rect 225234 82894 225854 118338
rect 225234 82658 225266 82894
rect 225502 82658 225586 82894
rect 225822 82658 225854 82894
rect 225234 82574 225854 82658
rect 225234 82338 225266 82574
rect 225502 82338 225586 82574
rect 225822 82338 225854 82574
rect 225234 46894 225854 82338
rect 225234 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 225854 46894
rect 225234 46574 225854 46658
rect 225234 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 225854 46574
rect 225234 10894 225854 46338
rect 225234 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 225854 10894
rect 225234 10574 225854 10658
rect 225234 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 225854 10574
rect 225234 -4186 225854 10338
rect 225234 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 225854 -4186
rect 225234 -4506 225854 -4422
rect 225234 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 225854 -4506
rect 225234 -5734 225854 -4742
rect 228954 698614 229574 710042
rect 246954 711558 247574 711590
rect 246954 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 247574 711558
rect 246954 711238 247574 711322
rect 246954 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 247574 711238
rect 243234 709638 243854 709670
rect 243234 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 243854 709638
rect 243234 709318 243854 709402
rect 243234 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 243854 709318
rect 239514 707718 240134 707750
rect 239514 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 240134 707718
rect 239514 707398 240134 707482
rect 239514 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 240134 707398
rect 235794 705798 236414 705830
rect 235794 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 236414 705798
rect 235794 705478 236414 705562
rect 235794 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 236414 705478
rect 235211 700500 235277 700501
rect 235211 700436 235212 700500
rect 235276 700436 235277 700500
rect 235211 700435 235277 700436
rect 228954 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 229574 698614
rect 228954 698294 229574 698378
rect 228954 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 229574 698294
rect 228954 662614 229574 698058
rect 228954 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 229574 662614
rect 228954 662294 229574 662378
rect 228954 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 229574 662294
rect 228954 626614 229574 662058
rect 228954 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 229574 626614
rect 228954 626294 229574 626378
rect 228954 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 229574 626294
rect 228954 590614 229574 626058
rect 228954 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 229574 590614
rect 228954 590294 229574 590378
rect 228954 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 229574 590294
rect 228954 554614 229574 590058
rect 228954 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 229574 554614
rect 228954 554294 229574 554378
rect 228954 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 229574 554294
rect 228954 518614 229574 554058
rect 228954 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 229574 518614
rect 228954 518294 229574 518378
rect 228954 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 229574 518294
rect 228954 482614 229574 518058
rect 228954 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 229574 482614
rect 228954 482294 229574 482378
rect 228954 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 229574 482294
rect 228954 446614 229574 482058
rect 228954 446378 228986 446614
rect 229222 446378 229306 446614
rect 229542 446378 229574 446614
rect 228954 446294 229574 446378
rect 228954 446058 228986 446294
rect 229222 446058 229306 446294
rect 229542 446058 229574 446294
rect 228954 410614 229574 446058
rect 228954 410378 228986 410614
rect 229222 410378 229306 410614
rect 229542 410378 229574 410614
rect 228954 410294 229574 410378
rect 228954 410058 228986 410294
rect 229222 410058 229306 410294
rect 229542 410058 229574 410294
rect 228954 374614 229574 410058
rect 228954 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 229574 374614
rect 228954 374294 229574 374378
rect 228954 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 229574 374294
rect 228954 338614 229574 374058
rect 228954 338378 228986 338614
rect 229222 338378 229306 338614
rect 229542 338378 229574 338614
rect 228954 338294 229574 338378
rect 228954 338058 228986 338294
rect 229222 338058 229306 338294
rect 229542 338058 229574 338294
rect 228954 302614 229574 338058
rect 228954 302378 228986 302614
rect 229222 302378 229306 302614
rect 229542 302378 229574 302614
rect 228954 302294 229574 302378
rect 228954 302058 228986 302294
rect 229222 302058 229306 302294
rect 229542 302058 229574 302294
rect 228954 266614 229574 302058
rect 228954 266378 228986 266614
rect 229222 266378 229306 266614
rect 229542 266378 229574 266614
rect 228954 266294 229574 266378
rect 228954 266058 228986 266294
rect 229222 266058 229306 266294
rect 229542 266058 229574 266294
rect 228954 230614 229574 266058
rect 228954 230378 228986 230614
rect 229222 230378 229306 230614
rect 229542 230378 229574 230614
rect 228954 230294 229574 230378
rect 228954 230058 228986 230294
rect 229222 230058 229306 230294
rect 229542 230058 229574 230294
rect 228954 194614 229574 230058
rect 228954 194378 228986 194614
rect 229222 194378 229306 194614
rect 229542 194378 229574 194614
rect 228954 194294 229574 194378
rect 228954 194058 228986 194294
rect 229222 194058 229306 194294
rect 229542 194058 229574 194294
rect 228954 158614 229574 194058
rect 235214 176493 235274 700435
rect 235794 669454 236414 705242
rect 237971 700636 238037 700637
rect 237971 700572 237972 700636
rect 238036 700572 238037 700636
rect 237971 700571 238037 700572
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235395 618356 235461 618357
rect 235395 618292 235396 618356
rect 235460 618292 235461 618356
rect 235395 618291 235461 618292
rect 235398 176629 235458 618291
rect 235794 597454 236414 632898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 561454 236414 596898
rect 235794 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 236414 561454
rect 235794 561134 236414 561218
rect 235794 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 236414 561134
rect 235794 525454 236414 560898
rect 235794 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 236414 525454
rect 235794 525134 236414 525218
rect 235794 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 236414 525134
rect 235794 489454 236414 524898
rect 235794 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 236414 489454
rect 235794 489134 236414 489218
rect 235794 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 236414 489134
rect 235794 453454 236414 488898
rect 235794 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 236414 453454
rect 235794 453134 236414 453218
rect 235794 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 236414 453134
rect 235794 417454 236414 452898
rect 235794 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 236414 417454
rect 235794 417134 236414 417218
rect 235794 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 236414 417134
rect 235794 381454 236414 416898
rect 235794 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 236414 381454
rect 235794 381134 236414 381218
rect 235794 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 236414 381134
rect 235794 345454 236414 380898
rect 235794 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 236414 345454
rect 235794 345134 236414 345218
rect 235794 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 236414 345134
rect 235794 309454 236414 344898
rect 235794 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 236414 309454
rect 235794 309134 236414 309218
rect 235794 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 236414 309134
rect 235794 273454 236414 308898
rect 235794 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 236414 273454
rect 235794 273134 236414 273218
rect 235794 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 236414 273134
rect 235794 237454 236414 272898
rect 235794 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 236414 237454
rect 235794 237134 236414 237218
rect 235794 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 236414 237134
rect 235794 201454 236414 236898
rect 235794 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 236414 201454
rect 235794 201134 236414 201218
rect 235794 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 236414 201134
rect 235395 176628 235461 176629
rect 235395 176564 235396 176628
rect 235460 176564 235461 176628
rect 235395 176563 235461 176564
rect 235211 176492 235277 176493
rect 235211 176428 235212 176492
rect 235276 176428 235277 176492
rect 235211 176427 235277 176428
rect 228954 158378 228986 158614
rect 229222 158378 229306 158614
rect 229542 158378 229574 158614
rect 228954 158294 229574 158378
rect 228954 158058 228986 158294
rect 229222 158058 229306 158294
rect 229542 158058 229574 158294
rect 228954 122614 229574 158058
rect 228954 122378 228986 122614
rect 229222 122378 229306 122614
rect 229542 122378 229574 122614
rect 228954 122294 229574 122378
rect 228954 122058 228986 122294
rect 229222 122058 229306 122294
rect 229542 122058 229574 122294
rect 228954 86614 229574 122058
rect 228954 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 229574 86614
rect 228954 86294 229574 86378
rect 228954 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 229574 86294
rect 228954 50614 229574 86058
rect 228954 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 229574 50614
rect 228954 50294 229574 50378
rect 228954 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 229574 50294
rect 228954 14614 229574 50058
rect 228954 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 229574 14614
rect 228954 14294 229574 14378
rect 228954 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 229574 14294
rect 210954 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 211574 -7066
rect 210954 -7386 211574 -7302
rect 210954 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 211574 -7386
rect 210954 -7654 211574 -7622
rect 228954 -6106 229574 14058
rect 235794 165454 236414 200898
rect 237974 179621 238034 700571
rect 239259 700364 239325 700365
rect 239259 700300 239260 700364
rect 239324 700300 239325 700364
rect 239259 700299 239325 700300
rect 238155 456924 238221 456925
rect 238155 456860 238156 456924
rect 238220 456860 238221 456924
rect 238155 456859 238221 456860
rect 238158 377909 238218 456859
rect 238339 451484 238405 451485
rect 238339 451420 238340 451484
rect 238404 451420 238405 451484
rect 238339 451419 238405 451420
rect 238342 379269 238402 451419
rect 238339 379268 238405 379269
rect 238339 379204 238340 379268
rect 238404 379204 238405 379268
rect 238339 379203 238405 379204
rect 238155 377908 238221 377909
rect 238155 377844 238156 377908
rect 238220 377844 238221 377908
rect 238155 377843 238221 377844
rect 238155 277676 238221 277677
rect 238155 277612 238156 277676
rect 238220 277612 238221 277676
rect 238155 277611 238221 277612
rect 238158 198525 238218 277611
rect 238339 268564 238405 268565
rect 238339 268500 238340 268564
rect 238404 268500 238405 268564
rect 238339 268499 238405 268500
rect 238342 200837 238402 268499
rect 238523 262444 238589 262445
rect 238523 262380 238524 262444
rect 238588 262380 238589 262444
rect 238523 262379 238589 262380
rect 238339 200836 238405 200837
rect 238339 200772 238340 200836
rect 238404 200772 238405 200836
rect 238339 200771 238405 200772
rect 238155 198524 238221 198525
rect 238155 198460 238156 198524
rect 238220 198460 238221 198524
rect 238155 198459 238221 198460
rect 238526 197573 238586 262379
rect 238523 197572 238589 197573
rect 238523 197508 238524 197572
rect 238588 197508 238589 197572
rect 238523 197507 238589 197508
rect 237971 179620 238037 179621
rect 237971 179556 237972 179620
rect 238036 179556 238037 179620
rect 237971 179555 238037 179556
rect 239262 178941 239322 700299
rect 239514 673174 240134 707162
rect 239514 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 240134 673174
rect 239514 672854 240134 672938
rect 239514 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 240134 672854
rect 239514 637174 240134 672618
rect 239514 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 240134 637174
rect 239514 636854 240134 636938
rect 239514 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 240134 636854
rect 239514 601174 240134 636618
rect 239514 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 240134 601174
rect 239514 600854 240134 600938
rect 239514 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 240134 600854
rect 239514 565174 240134 600618
rect 239514 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 240134 565174
rect 239514 564854 240134 564938
rect 239514 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 240134 564854
rect 239514 529174 240134 564618
rect 239514 528938 239546 529174
rect 239782 528938 239866 529174
rect 240102 528938 240134 529174
rect 239514 528854 240134 528938
rect 239514 528618 239546 528854
rect 239782 528618 239866 528854
rect 240102 528618 240134 528854
rect 239514 493174 240134 528618
rect 239514 492938 239546 493174
rect 239782 492938 239866 493174
rect 240102 492938 240134 493174
rect 239514 492854 240134 492938
rect 239514 492618 239546 492854
rect 239782 492618 239866 492854
rect 240102 492618 240134 492854
rect 239514 482000 240134 492618
rect 243234 676894 243854 709082
rect 243234 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 243854 676894
rect 243234 676574 243854 676658
rect 243234 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 243854 676574
rect 243234 640894 243854 676338
rect 243234 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 243854 640894
rect 243234 640574 243854 640658
rect 243234 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 243854 640574
rect 243234 604894 243854 640338
rect 243234 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 243854 604894
rect 243234 604574 243854 604658
rect 243234 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 243854 604574
rect 243234 568894 243854 604338
rect 243234 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 243854 568894
rect 243234 568574 243854 568658
rect 243234 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 243854 568574
rect 243234 532894 243854 568338
rect 243234 532658 243266 532894
rect 243502 532658 243586 532894
rect 243822 532658 243854 532894
rect 243234 532574 243854 532658
rect 243234 532338 243266 532574
rect 243502 532338 243586 532574
rect 243822 532338 243854 532574
rect 243234 496894 243854 532338
rect 243234 496658 243266 496894
rect 243502 496658 243586 496894
rect 243822 496658 243854 496894
rect 243234 496574 243854 496658
rect 243234 496338 243266 496574
rect 243502 496338 243586 496574
rect 243822 496338 243854 496574
rect 243234 482000 243854 496338
rect 246954 680614 247574 711002
rect 264954 710598 265574 711590
rect 264954 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 265574 710598
rect 264954 710278 265574 710362
rect 264954 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 265574 710278
rect 261234 708678 261854 709670
rect 261234 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 261854 708678
rect 261234 708358 261854 708442
rect 261234 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 261854 708358
rect 257514 706758 258134 707750
rect 257514 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 258134 706758
rect 257514 706438 258134 706522
rect 257514 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 258134 706438
rect 246954 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 247574 680614
rect 246954 680294 247574 680378
rect 246954 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 247574 680294
rect 246954 644614 247574 680058
rect 246954 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 247574 644614
rect 246954 644294 247574 644378
rect 246954 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 247574 644294
rect 246954 608614 247574 644058
rect 246954 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 247574 608614
rect 246954 608294 247574 608378
rect 246954 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 247574 608294
rect 246954 572614 247574 608058
rect 246954 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 247574 572614
rect 246954 572294 247574 572378
rect 246954 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 247574 572294
rect 246954 536614 247574 572058
rect 246954 536378 246986 536614
rect 247222 536378 247306 536614
rect 247542 536378 247574 536614
rect 246954 536294 247574 536378
rect 246954 536058 246986 536294
rect 247222 536058 247306 536294
rect 247542 536058 247574 536294
rect 246954 500614 247574 536058
rect 246954 500378 246986 500614
rect 247222 500378 247306 500614
rect 247542 500378 247574 500614
rect 246954 500294 247574 500378
rect 246954 500058 246986 500294
rect 247222 500058 247306 500294
rect 247542 500058 247574 500294
rect 246954 482000 247574 500058
rect 253794 704838 254414 705830
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 543454 254414 578898
rect 253794 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 254414 543454
rect 253794 543134 254414 543218
rect 253794 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 254414 543134
rect 253794 507454 254414 542898
rect 253794 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 254414 507454
rect 253794 507134 254414 507218
rect 253794 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 254414 507134
rect 253794 482000 254414 506898
rect 257514 691174 258134 706202
rect 257514 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 258134 691174
rect 257514 690854 258134 690938
rect 257514 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 258134 690854
rect 257514 655174 258134 690618
rect 257514 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 258134 655174
rect 257514 654854 258134 654938
rect 257514 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 258134 654854
rect 257514 619174 258134 654618
rect 257514 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 258134 619174
rect 257514 618854 258134 618938
rect 257514 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 258134 618854
rect 257514 583174 258134 618618
rect 257514 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 258134 583174
rect 257514 582854 258134 582938
rect 257514 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 258134 582854
rect 257514 547174 258134 582618
rect 257514 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 258134 547174
rect 257514 546854 258134 546938
rect 257514 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 258134 546854
rect 257514 511174 258134 546618
rect 257514 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 258134 511174
rect 257514 510854 258134 510938
rect 257514 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 258134 510854
rect 257514 482000 258134 510618
rect 261234 694894 261854 708122
rect 261234 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 261854 694894
rect 261234 694574 261854 694658
rect 261234 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 261854 694574
rect 261234 658894 261854 694338
rect 261234 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 261854 658894
rect 261234 658574 261854 658658
rect 261234 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 261854 658574
rect 261234 622894 261854 658338
rect 261234 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 261854 622894
rect 261234 622574 261854 622658
rect 261234 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 261854 622574
rect 261234 586894 261854 622338
rect 261234 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 261854 586894
rect 261234 586574 261854 586658
rect 261234 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 261854 586574
rect 261234 550894 261854 586338
rect 261234 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 261854 550894
rect 261234 550574 261854 550658
rect 261234 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 261854 550574
rect 261234 514894 261854 550338
rect 261234 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 261854 514894
rect 261234 514574 261854 514658
rect 261234 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 261854 514574
rect 261234 482000 261854 514338
rect 264954 698614 265574 710042
rect 282954 711558 283574 711590
rect 282954 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 283574 711558
rect 282954 711238 283574 711322
rect 282954 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 283574 711238
rect 279234 709638 279854 709670
rect 279234 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 279854 709638
rect 279234 709318 279854 709402
rect 279234 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 279854 709318
rect 275514 707718 276134 707750
rect 275514 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 276134 707718
rect 275514 707398 276134 707482
rect 275514 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 276134 707398
rect 264954 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 265574 698614
rect 264954 698294 265574 698378
rect 264954 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 265574 698294
rect 264954 662614 265574 698058
rect 264954 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 265574 662614
rect 264954 662294 265574 662378
rect 264954 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 265574 662294
rect 264954 626614 265574 662058
rect 264954 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 265574 626614
rect 264954 626294 265574 626378
rect 264954 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 265574 626294
rect 264954 590614 265574 626058
rect 264954 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 265574 590614
rect 264954 590294 265574 590378
rect 264954 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 265574 590294
rect 264954 554614 265574 590058
rect 264954 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 265574 554614
rect 264954 554294 265574 554378
rect 264954 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 265574 554294
rect 264954 518614 265574 554058
rect 264954 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 265574 518614
rect 264954 518294 265574 518378
rect 264954 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 265574 518294
rect 264954 482614 265574 518058
rect 264954 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 265574 482614
rect 264954 482294 265574 482378
rect 264954 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 265574 482294
rect 264954 482000 265574 482058
rect 271794 705798 272414 705830
rect 271794 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 272414 705798
rect 271794 705478 272414 705562
rect 271794 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 272414 705478
rect 271794 669454 272414 705242
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 561454 272414 596898
rect 271794 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 272414 561454
rect 271794 561134 272414 561218
rect 271794 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 272414 561134
rect 271794 525454 272414 560898
rect 271794 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 272414 525454
rect 271794 525134 272414 525218
rect 271794 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 272414 525134
rect 271794 489454 272414 524898
rect 271794 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 272414 489454
rect 271794 489134 272414 489218
rect 271794 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 272414 489134
rect 271794 482000 272414 488898
rect 275514 673174 276134 707162
rect 275514 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 276134 673174
rect 275514 672854 276134 672938
rect 275514 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 276134 672854
rect 275514 637174 276134 672618
rect 275514 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 276134 637174
rect 275514 636854 276134 636938
rect 275514 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 276134 636854
rect 275514 601174 276134 636618
rect 275514 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 276134 601174
rect 275514 600854 276134 600938
rect 275514 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 276134 600854
rect 275514 565174 276134 600618
rect 275514 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 276134 565174
rect 275514 564854 276134 564938
rect 275514 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 276134 564854
rect 275514 529174 276134 564618
rect 275514 528938 275546 529174
rect 275782 528938 275866 529174
rect 276102 528938 276134 529174
rect 275514 528854 276134 528938
rect 275514 528618 275546 528854
rect 275782 528618 275866 528854
rect 276102 528618 276134 528854
rect 275514 493174 276134 528618
rect 275514 492938 275546 493174
rect 275782 492938 275866 493174
rect 276102 492938 276134 493174
rect 275514 492854 276134 492938
rect 275514 492618 275546 492854
rect 275782 492618 275866 492854
rect 276102 492618 276134 492854
rect 275514 482000 276134 492618
rect 279234 676894 279854 709082
rect 279234 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 279854 676894
rect 279234 676574 279854 676658
rect 279234 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 279854 676574
rect 279234 640894 279854 676338
rect 279234 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 279854 640894
rect 279234 640574 279854 640658
rect 279234 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 279854 640574
rect 279234 604894 279854 640338
rect 279234 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 279854 604894
rect 279234 604574 279854 604658
rect 279234 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 279854 604574
rect 279234 568894 279854 604338
rect 279234 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 279854 568894
rect 279234 568574 279854 568658
rect 279234 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 279854 568574
rect 279234 532894 279854 568338
rect 279234 532658 279266 532894
rect 279502 532658 279586 532894
rect 279822 532658 279854 532894
rect 279234 532574 279854 532658
rect 279234 532338 279266 532574
rect 279502 532338 279586 532574
rect 279822 532338 279854 532574
rect 279234 496894 279854 532338
rect 279234 496658 279266 496894
rect 279502 496658 279586 496894
rect 279822 496658 279854 496894
rect 279234 496574 279854 496658
rect 279234 496338 279266 496574
rect 279502 496338 279586 496574
rect 279822 496338 279854 496574
rect 279234 482000 279854 496338
rect 282954 680614 283574 711002
rect 300954 710598 301574 711590
rect 300954 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 301574 710598
rect 300954 710278 301574 710362
rect 300954 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 301574 710278
rect 297234 708678 297854 709670
rect 297234 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 297854 708678
rect 297234 708358 297854 708442
rect 297234 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 297854 708358
rect 293514 706758 294134 707750
rect 293514 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 294134 706758
rect 293514 706438 294134 706522
rect 293514 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 294134 706438
rect 282954 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 283574 680614
rect 282954 680294 283574 680378
rect 282954 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 283574 680294
rect 282954 644614 283574 680058
rect 282954 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 283574 644614
rect 282954 644294 283574 644378
rect 282954 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 283574 644294
rect 282954 608614 283574 644058
rect 282954 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 283574 608614
rect 282954 608294 283574 608378
rect 282954 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 283574 608294
rect 282954 572614 283574 608058
rect 282954 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 283574 572614
rect 282954 572294 283574 572378
rect 282954 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 283574 572294
rect 282954 536614 283574 572058
rect 282954 536378 282986 536614
rect 283222 536378 283306 536614
rect 283542 536378 283574 536614
rect 282954 536294 283574 536378
rect 282954 536058 282986 536294
rect 283222 536058 283306 536294
rect 283542 536058 283574 536294
rect 282954 500614 283574 536058
rect 282954 500378 282986 500614
rect 283222 500378 283306 500614
rect 283542 500378 283574 500614
rect 282954 500294 283574 500378
rect 282954 500058 282986 500294
rect 283222 500058 283306 500294
rect 283542 500058 283574 500294
rect 282954 482000 283574 500058
rect 289794 704838 290414 705830
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 543454 290414 578898
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289794 507454 290414 542898
rect 289794 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 290414 507454
rect 289794 507134 290414 507218
rect 289794 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 290414 507134
rect 289794 482000 290414 506898
rect 293514 691174 294134 706202
rect 293514 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 294134 691174
rect 293514 690854 294134 690938
rect 293514 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 294134 690854
rect 293514 655174 294134 690618
rect 293514 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 294134 655174
rect 293514 654854 294134 654938
rect 293514 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 294134 654854
rect 293514 619174 294134 654618
rect 293514 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 294134 619174
rect 293514 618854 294134 618938
rect 293514 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 294134 618854
rect 293514 583174 294134 618618
rect 293514 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 294134 583174
rect 293514 582854 294134 582938
rect 293514 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 294134 582854
rect 293514 547174 294134 582618
rect 293514 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 294134 547174
rect 293514 546854 294134 546938
rect 293514 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 294134 546854
rect 293514 511174 294134 546618
rect 293514 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 294134 511174
rect 293514 510854 294134 510938
rect 293514 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 294134 510854
rect 293514 482000 294134 510618
rect 297234 694894 297854 708122
rect 297234 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 297854 694894
rect 297234 694574 297854 694658
rect 297234 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 297854 694574
rect 297234 658894 297854 694338
rect 297234 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 297854 658894
rect 297234 658574 297854 658658
rect 297234 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 297854 658574
rect 297234 622894 297854 658338
rect 297234 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 297854 622894
rect 297234 622574 297854 622658
rect 297234 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 297854 622574
rect 297234 586894 297854 622338
rect 297234 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 297854 586894
rect 297234 586574 297854 586658
rect 297234 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 297854 586574
rect 297234 550894 297854 586338
rect 297234 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 297854 550894
rect 297234 550574 297854 550658
rect 297234 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 297854 550574
rect 297234 514894 297854 550338
rect 297234 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 297854 514894
rect 297234 514574 297854 514658
rect 297234 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 297854 514574
rect 297234 482000 297854 514338
rect 300954 698614 301574 710042
rect 318954 711558 319574 711590
rect 318954 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 319574 711558
rect 318954 711238 319574 711322
rect 318954 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 319574 711238
rect 315234 709638 315854 709670
rect 315234 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 315854 709638
rect 315234 709318 315854 709402
rect 315234 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 315854 709318
rect 311514 707718 312134 707750
rect 311514 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 312134 707718
rect 311514 707398 312134 707482
rect 311514 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 312134 707398
rect 300954 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 301574 698614
rect 300954 698294 301574 698378
rect 300954 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 301574 698294
rect 300954 662614 301574 698058
rect 300954 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 301574 662614
rect 300954 662294 301574 662378
rect 300954 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 301574 662294
rect 300954 626614 301574 662058
rect 300954 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 301574 626614
rect 300954 626294 301574 626378
rect 300954 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 301574 626294
rect 300954 590614 301574 626058
rect 300954 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 301574 590614
rect 300954 590294 301574 590378
rect 300954 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 301574 590294
rect 300954 554614 301574 590058
rect 300954 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 301574 554614
rect 300954 554294 301574 554378
rect 300954 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 301574 554294
rect 300954 518614 301574 554058
rect 300954 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 301574 518614
rect 300954 518294 301574 518378
rect 300954 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 301574 518294
rect 300954 482614 301574 518058
rect 300954 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 301574 482614
rect 300954 482294 301574 482378
rect 300954 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 301574 482294
rect 300954 482000 301574 482058
rect 307794 705798 308414 705830
rect 307794 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 308414 705798
rect 307794 705478 308414 705562
rect 307794 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 308414 705478
rect 307794 669454 308414 705242
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 561454 308414 596898
rect 307794 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 308414 561454
rect 307794 561134 308414 561218
rect 307794 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 308414 561134
rect 307794 525454 308414 560898
rect 307794 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 308414 525454
rect 307794 525134 308414 525218
rect 307794 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 308414 525134
rect 307794 489454 308414 524898
rect 307794 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 308414 489454
rect 307794 489134 308414 489218
rect 307794 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 308414 489134
rect 307794 482000 308414 488898
rect 311514 673174 312134 707162
rect 311514 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 312134 673174
rect 311514 672854 312134 672938
rect 311514 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 312134 672854
rect 311514 637174 312134 672618
rect 311514 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 312134 637174
rect 311514 636854 312134 636938
rect 311514 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 312134 636854
rect 311514 601174 312134 636618
rect 311514 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 312134 601174
rect 311514 600854 312134 600938
rect 311514 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 312134 600854
rect 311514 565174 312134 600618
rect 311514 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 312134 565174
rect 311514 564854 312134 564938
rect 311514 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 312134 564854
rect 311514 529174 312134 564618
rect 311514 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 312134 529174
rect 311514 528854 312134 528938
rect 311514 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 312134 528854
rect 311514 493174 312134 528618
rect 311514 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 312134 493174
rect 311514 492854 312134 492938
rect 311514 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 312134 492854
rect 311514 482000 312134 492618
rect 315234 676894 315854 709082
rect 315234 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 315854 676894
rect 315234 676574 315854 676658
rect 315234 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 315854 676574
rect 315234 640894 315854 676338
rect 315234 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 315854 640894
rect 315234 640574 315854 640658
rect 315234 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 315854 640574
rect 315234 604894 315854 640338
rect 315234 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 315854 604894
rect 315234 604574 315854 604658
rect 315234 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 315854 604574
rect 315234 568894 315854 604338
rect 315234 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 315854 568894
rect 315234 568574 315854 568658
rect 315234 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 315854 568574
rect 315234 532894 315854 568338
rect 315234 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 315854 532894
rect 315234 532574 315854 532658
rect 315234 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 315854 532574
rect 315234 496894 315854 532338
rect 315234 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 315854 496894
rect 315234 496574 315854 496658
rect 315234 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 315854 496574
rect 315234 482000 315854 496338
rect 318954 680614 319574 711002
rect 336954 710598 337574 711590
rect 336954 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 337574 710598
rect 336954 710278 337574 710362
rect 336954 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 337574 710278
rect 333234 708678 333854 709670
rect 333234 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 333854 708678
rect 333234 708358 333854 708442
rect 333234 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 333854 708358
rect 329514 706758 330134 707750
rect 329514 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 330134 706758
rect 329514 706438 330134 706522
rect 329514 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 330134 706438
rect 318954 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 319574 680614
rect 318954 680294 319574 680378
rect 318954 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 319574 680294
rect 318954 644614 319574 680058
rect 318954 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 319574 644614
rect 318954 644294 319574 644378
rect 318954 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 319574 644294
rect 318954 608614 319574 644058
rect 318954 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 319574 608614
rect 318954 608294 319574 608378
rect 318954 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 319574 608294
rect 318954 572614 319574 608058
rect 318954 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 319574 572614
rect 318954 572294 319574 572378
rect 318954 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 319574 572294
rect 318954 536614 319574 572058
rect 318954 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 319574 536614
rect 318954 536294 319574 536378
rect 318954 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 319574 536294
rect 318954 500614 319574 536058
rect 318954 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 319574 500614
rect 318954 500294 319574 500378
rect 318954 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 319574 500294
rect 318954 482000 319574 500058
rect 325794 704838 326414 705830
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 543454 326414 578898
rect 325794 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 326414 543454
rect 325794 543134 326414 543218
rect 325794 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 326414 543134
rect 325794 507454 326414 542898
rect 325794 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 326414 507454
rect 325794 507134 326414 507218
rect 325794 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 326414 507134
rect 325794 482000 326414 506898
rect 329514 691174 330134 706202
rect 329514 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 330134 691174
rect 329514 690854 330134 690938
rect 329514 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 330134 690854
rect 329514 655174 330134 690618
rect 329514 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 330134 655174
rect 329514 654854 330134 654938
rect 329514 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 330134 654854
rect 329514 619174 330134 654618
rect 329514 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 330134 619174
rect 329514 618854 330134 618938
rect 329514 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 330134 618854
rect 329514 583174 330134 618618
rect 329514 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 330134 583174
rect 329514 582854 330134 582938
rect 329514 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 330134 582854
rect 329514 547174 330134 582618
rect 329514 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 330134 547174
rect 329514 546854 330134 546938
rect 329514 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 330134 546854
rect 329514 511174 330134 546618
rect 329514 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 330134 511174
rect 329514 510854 330134 510938
rect 329514 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 330134 510854
rect 329514 482000 330134 510618
rect 333234 694894 333854 708122
rect 333234 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 333854 694894
rect 333234 694574 333854 694658
rect 333234 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 333854 694574
rect 333234 658894 333854 694338
rect 333234 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 333854 658894
rect 333234 658574 333854 658658
rect 333234 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 333854 658574
rect 333234 622894 333854 658338
rect 333234 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 333854 622894
rect 333234 622574 333854 622658
rect 333234 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 333854 622574
rect 333234 586894 333854 622338
rect 333234 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 333854 586894
rect 333234 586574 333854 586658
rect 333234 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 333854 586574
rect 333234 550894 333854 586338
rect 333234 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 333854 550894
rect 333234 550574 333854 550658
rect 333234 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 333854 550574
rect 333234 514894 333854 550338
rect 333234 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 333854 514894
rect 333234 514574 333854 514658
rect 333234 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 333854 514574
rect 333234 482000 333854 514338
rect 336954 698614 337574 710042
rect 354954 711558 355574 711590
rect 354954 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 355574 711558
rect 354954 711238 355574 711322
rect 354954 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 355574 711238
rect 351234 709638 351854 709670
rect 351234 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 351854 709638
rect 351234 709318 351854 709402
rect 351234 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 351854 709318
rect 347514 707718 348134 707750
rect 347514 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 348134 707718
rect 347514 707398 348134 707482
rect 347514 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 348134 707398
rect 336954 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 337574 698614
rect 336954 698294 337574 698378
rect 336954 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 337574 698294
rect 336954 662614 337574 698058
rect 336954 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 337574 662614
rect 336954 662294 337574 662378
rect 336954 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 337574 662294
rect 336954 626614 337574 662058
rect 336954 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 337574 626614
rect 336954 626294 337574 626378
rect 336954 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 337574 626294
rect 336954 590614 337574 626058
rect 336954 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 337574 590614
rect 336954 590294 337574 590378
rect 336954 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 337574 590294
rect 336954 554614 337574 590058
rect 336954 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 337574 554614
rect 336954 554294 337574 554378
rect 336954 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 337574 554294
rect 336954 518614 337574 554058
rect 336954 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 337574 518614
rect 336954 518294 337574 518378
rect 336954 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 337574 518294
rect 336954 482614 337574 518058
rect 336954 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 337574 482614
rect 336954 482294 337574 482378
rect 336954 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 337574 482294
rect 336954 482000 337574 482058
rect 343794 705798 344414 705830
rect 343794 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 344414 705798
rect 343794 705478 344414 705562
rect 343794 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 344414 705478
rect 343794 669454 344414 705242
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 561454 344414 596898
rect 343794 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 344414 561454
rect 343794 561134 344414 561218
rect 343794 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 344414 561134
rect 343794 525454 344414 560898
rect 343794 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 344414 525454
rect 343794 525134 344414 525218
rect 343794 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 344414 525134
rect 343794 489454 344414 524898
rect 343794 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 344414 489454
rect 343794 489134 344414 489218
rect 343794 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 344414 489134
rect 343794 482000 344414 488898
rect 347514 673174 348134 707162
rect 347514 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 348134 673174
rect 347514 672854 348134 672938
rect 347514 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 348134 672854
rect 347514 637174 348134 672618
rect 347514 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 348134 637174
rect 347514 636854 348134 636938
rect 347514 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 348134 636854
rect 347514 601174 348134 636618
rect 347514 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 348134 601174
rect 347514 600854 348134 600938
rect 347514 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 348134 600854
rect 347514 565174 348134 600618
rect 347514 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 348134 565174
rect 347514 564854 348134 564938
rect 347514 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 348134 564854
rect 347514 529174 348134 564618
rect 347514 528938 347546 529174
rect 347782 528938 347866 529174
rect 348102 528938 348134 529174
rect 347514 528854 348134 528938
rect 347514 528618 347546 528854
rect 347782 528618 347866 528854
rect 348102 528618 348134 528854
rect 347514 493174 348134 528618
rect 347514 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 348134 493174
rect 347514 492854 348134 492938
rect 347514 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 348134 492854
rect 347514 482000 348134 492618
rect 351234 676894 351854 709082
rect 351234 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 351854 676894
rect 351234 676574 351854 676658
rect 351234 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 351854 676574
rect 351234 640894 351854 676338
rect 351234 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 351854 640894
rect 351234 640574 351854 640658
rect 351234 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 351854 640574
rect 351234 604894 351854 640338
rect 351234 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 351854 604894
rect 351234 604574 351854 604658
rect 351234 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 351854 604574
rect 351234 568894 351854 604338
rect 351234 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 351854 568894
rect 351234 568574 351854 568658
rect 351234 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 351854 568574
rect 351234 532894 351854 568338
rect 351234 532658 351266 532894
rect 351502 532658 351586 532894
rect 351822 532658 351854 532894
rect 351234 532574 351854 532658
rect 351234 532338 351266 532574
rect 351502 532338 351586 532574
rect 351822 532338 351854 532574
rect 351234 496894 351854 532338
rect 351234 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 351854 496894
rect 351234 496574 351854 496658
rect 351234 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 351854 496574
rect 351234 482000 351854 496338
rect 354954 680614 355574 711002
rect 372954 710598 373574 711590
rect 372954 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 373574 710598
rect 372954 710278 373574 710362
rect 372954 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 373574 710278
rect 369234 708678 369854 709670
rect 369234 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 369854 708678
rect 369234 708358 369854 708442
rect 369234 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 369854 708358
rect 365514 706758 366134 707750
rect 365514 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 366134 706758
rect 365514 706438 366134 706522
rect 365514 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 366134 706438
rect 354954 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 355574 680614
rect 354954 680294 355574 680378
rect 354954 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 355574 680294
rect 354954 644614 355574 680058
rect 354954 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 355574 644614
rect 354954 644294 355574 644378
rect 354954 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 355574 644294
rect 354954 608614 355574 644058
rect 354954 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 355574 608614
rect 354954 608294 355574 608378
rect 354954 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 355574 608294
rect 354954 572614 355574 608058
rect 354954 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 355574 572614
rect 354954 572294 355574 572378
rect 354954 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 355574 572294
rect 354954 536614 355574 572058
rect 354954 536378 354986 536614
rect 355222 536378 355306 536614
rect 355542 536378 355574 536614
rect 354954 536294 355574 536378
rect 354954 536058 354986 536294
rect 355222 536058 355306 536294
rect 355542 536058 355574 536294
rect 354954 500614 355574 536058
rect 354954 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 355574 500614
rect 354954 500294 355574 500378
rect 354954 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 355574 500294
rect 354954 482000 355574 500058
rect 361794 704838 362414 705830
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 361794 482000 362414 506898
rect 365514 691174 366134 706202
rect 365514 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 366134 691174
rect 365514 690854 366134 690938
rect 365514 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 366134 690854
rect 365514 655174 366134 690618
rect 365514 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 366134 655174
rect 365514 654854 366134 654938
rect 365514 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 366134 654854
rect 365514 619174 366134 654618
rect 365514 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 366134 619174
rect 365514 618854 366134 618938
rect 365514 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 366134 618854
rect 365514 583174 366134 618618
rect 365514 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 366134 583174
rect 365514 582854 366134 582938
rect 365514 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 366134 582854
rect 365514 547174 366134 582618
rect 365514 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 366134 547174
rect 365514 546854 366134 546938
rect 365514 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 366134 546854
rect 365514 511174 366134 546618
rect 365514 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 366134 511174
rect 365514 510854 366134 510938
rect 365514 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 366134 510854
rect 365514 482000 366134 510618
rect 369234 694894 369854 708122
rect 369234 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 369854 694894
rect 369234 694574 369854 694658
rect 369234 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 369854 694574
rect 369234 658894 369854 694338
rect 369234 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 369854 658894
rect 369234 658574 369854 658658
rect 369234 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 369854 658574
rect 369234 622894 369854 658338
rect 369234 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 369854 622894
rect 369234 622574 369854 622658
rect 369234 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 369854 622574
rect 369234 586894 369854 622338
rect 369234 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 369854 586894
rect 369234 586574 369854 586658
rect 369234 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 369854 586574
rect 369234 550894 369854 586338
rect 369234 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 369854 550894
rect 369234 550574 369854 550658
rect 369234 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 369854 550574
rect 369234 514894 369854 550338
rect 369234 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 369854 514894
rect 369234 514574 369854 514658
rect 369234 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 369854 514574
rect 369234 482000 369854 514338
rect 372954 698614 373574 710042
rect 390954 711558 391574 711590
rect 390954 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 391574 711558
rect 390954 711238 391574 711322
rect 390954 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 391574 711238
rect 387234 709638 387854 709670
rect 387234 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 387854 709638
rect 387234 709318 387854 709402
rect 387234 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 387854 709318
rect 383514 707718 384134 707750
rect 383514 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 384134 707718
rect 383514 707398 384134 707482
rect 383514 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 384134 707398
rect 372954 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 373574 698614
rect 372954 698294 373574 698378
rect 372954 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 373574 698294
rect 372954 662614 373574 698058
rect 372954 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 373574 662614
rect 372954 662294 373574 662378
rect 372954 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 373574 662294
rect 372954 626614 373574 662058
rect 372954 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 373574 626614
rect 372954 626294 373574 626378
rect 372954 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 373574 626294
rect 372954 590614 373574 626058
rect 372954 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 373574 590614
rect 372954 590294 373574 590378
rect 372954 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 373574 590294
rect 372954 554614 373574 590058
rect 372954 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 373574 554614
rect 372954 554294 373574 554378
rect 372954 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 373574 554294
rect 372954 518614 373574 554058
rect 372954 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 373574 518614
rect 372954 518294 373574 518378
rect 372954 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 373574 518294
rect 372954 482614 373574 518058
rect 372954 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 373574 482614
rect 372954 482294 373574 482378
rect 372954 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 373574 482294
rect 372954 482000 373574 482058
rect 379794 705798 380414 705830
rect 379794 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 380414 705798
rect 379794 705478 380414 705562
rect 379794 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 380414 705478
rect 379794 669454 380414 705242
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 561454 380414 596898
rect 379794 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 380414 561454
rect 379794 561134 380414 561218
rect 379794 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 380414 561134
rect 379794 525454 380414 560898
rect 379794 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 380414 525454
rect 379794 525134 380414 525218
rect 379794 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 380414 525134
rect 379794 489454 380414 524898
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 379794 482000 380414 488898
rect 383514 673174 384134 707162
rect 383514 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 384134 673174
rect 383514 672854 384134 672938
rect 383514 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 384134 672854
rect 383514 637174 384134 672618
rect 383514 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 384134 637174
rect 383514 636854 384134 636938
rect 383514 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 384134 636854
rect 383514 601174 384134 636618
rect 383514 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 384134 601174
rect 383514 600854 384134 600938
rect 383514 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 384134 600854
rect 383514 565174 384134 600618
rect 383514 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 384134 565174
rect 383514 564854 384134 564938
rect 383514 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 384134 564854
rect 383514 529174 384134 564618
rect 383514 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 384134 529174
rect 383514 528854 384134 528938
rect 383514 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 384134 528854
rect 383514 493174 384134 528618
rect 383514 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 384134 493174
rect 383514 492854 384134 492938
rect 383514 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 384134 492854
rect 383514 482000 384134 492618
rect 387234 676894 387854 709082
rect 387234 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 387854 676894
rect 387234 676574 387854 676658
rect 387234 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 387854 676574
rect 387234 640894 387854 676338
rect 387234 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 387854 640894
rect 387234 640574 387854 640658
rect 387234 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 387854 640574
rect 387234 604894 387854 640338
rect 387234 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 387854 604894
rect 387234 604574 387854 604658
rect 387234 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 387854 604574
rect 387234 568894 387854 604338
rect 387234 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 387854 568894
rect 387234 568574 387854 568658
rect 387234 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 387854 568574
rect 387234 532894 387854 568338
rect 387234 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 387854 532894
rect 387234 532574 387854 532658
rect 387234 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 387854 532574
rect 387234 496894 387854 532338
rect 387234 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 387854 496894
rect 387234 496574 387854 496658
rect 387234 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 387854 496574
rect 387234 482000 387854 496338
rect 390954 680614 391574 711002
rect 408954 710598 409574 711590
rect 408954 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 409574 710598
rect 408954 710278 409574 710362
rect 408954 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 409574 710278
rect 405234 708678 405854 709670
rect 405234 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 405854 708678
rect 405234 708358 405854 708442
rect 405234 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 405854 708358
rect 401514 706758 402134 707750
rect 401514 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 402134 706758
rect 401514 706438 402134 706522
rect 401514 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 402134 706438
rect 390954 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 391574 680614
rect 390954 680294 391574 680378
rect 390954 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 391574 680294
rect 390954 644614 391574 680058
rect 390954 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 391574 644614
rect 390954 644294 391574 644378
rect 390954 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 391574 644294
rect 390954 608614 391574 644058
rect 390954 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 391574 608614
rect 390954 608294 391574 608378
rect 390954 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 391574 608294
rect 390954 572614 391574 608058
rect 390954 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 391574 572614
rect 390954 572294 391574 572378
rect 390954 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 391574 572294
rect 390954 536614 391574 572058
rect 390954 536378 390986 536614
rect 391222 536378 391306 536614
rect 391542 536378 391574 536614
rect 390954 536294 391574 536378
rect 390954 536058 390986 536294
rect 391222 536058 391306 536294
rect 391542 536058 391574 536294
rect 390954 500614 391574 536058
rect 390954 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 391574 500614
rect 390954 500294 391574 500378
rect 390954 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 391574 500294
rect 390954 482000 391574 500058
rect 397794 704838 398414 705830
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 482000 398414 506898
rect 401514 691174 402134 706202
rect 401514 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 402134 691174
rect 401514 690854 402134 690938
rect 401514 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 402134 690854
rect 401514 655174 402134 690618
rect 401514 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 402134 655174
rect 401514 654854 402134 654938
rect 401514 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 402134 654854
rect 401514 619174 402134 654618
rect 401514 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 402134 619174
rect 401514 618854 402134 618938
rect 401514 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 402134 618854
rect 401514 583174 402134 618618
rect 401514 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 402134 583174
rect 401514 582854 402134 582938
rect 401514 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 402134 582854
rect 401514 547174 402134 582618
rect 401514 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 402134 547174
rect 401514 546854 402134 546938
rect 401514 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 402134 546854
rect 401514 511174 402134 546618
rect 401514 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 402134 511174
rect 401514 510854 402134 510938
rect 401514 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 402134 510854
rect 401514 482000 402134 510618
rect 405234 694894 405854 708122
rect 405234 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 405854 694894
rect 405234 694574 405854 694658
rect 405234 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 405854 694574
rect 405234 658894 405854 694338
rect 405234 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 405854 658894
rect 405234 658574 405854 658658
rect 405234 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 405854 658574
rect 405234 622894 405854 658338
rect 405234 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 405854 622894
rect 405234 622574 405854 622658
rect 405234 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 405854 622574
rect 405234 586894 405854 622338
rect 405234 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 405854 586894
rect 405234 586574 405854 586658
rect 405234 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 405854 586574
rect 405234 550894 405854 586338
rect 405234 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 405854 550894
rect 405234 550574 405854 550658
rect 405234 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 405854 550574
rect 405234 514894 405854 550338
rect 405234 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 405854 514894
rect 405234 514574 405854 514658
rect 405234 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 405854 514574
rect 405234 482000 405854 514338
rect 408954 698614 409574 710042
rect 426954 711558 427574 711590
rect 426954 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 427574 711558
rect 426954 711238 427574 711322
rect 426954 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 427574 711238
rect 423234 709638 423854 709670
rect 423234 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 423854 709638
rect 423234 709318 423854 709402
rect 423234 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 423854 709318
rect 419514 707718 420134 707750
rect 419514 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 420134 707718
rect 419514 707398 420134 707482
rect 419514 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 420134 707398
rect 408954 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 409574 698614
rect 408954 698294 409574 698378
rect 408954 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 409574 698294
rect 408954 662614 409574 698058
rect 408954 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 409574 662614
rect 408954 662294 409574 662378
rect 408954 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 409574 662294
rect 408954 626614 409574 662058
rect 408954 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 409574 626614
rect 408954 626294 409574 626378
rect 408954 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 409574 626294
rect 408954 590614 409574 626058
rect 408954 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 409574 590614
rect 408954 590294 409574 590378
rect 408954 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 409574 590294
rect 408954 554614 409574 590058
rect 408954 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 409574 554614
rect 408954 554294 409574 554378
rect 408954 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 409574 554294
rect 408954 518614 409574 554058
rect 408954 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 409574 518614
rect 408954 518294 409574 518378
rect 408954 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 409574 518294
rect 408954 482614 409574 518058
rect 408954 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 409574 482614
rect 408954 482294 409574 482378
rect 408954 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 409574 482294
rect 408954 482000 409574 482058
rect 415794 705798 416414 705830
rect 415794 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 416414 705798
rect 415794 705478 416414 705562
rect 415794 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 416414 705478
rect 415794 669454 416414 705242
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 561454 416414 596898
rect 415794 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 416414 561454
rect 415794 561134 416414 561218
rect 415794 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 416414 561134
rect 415794 525454 416414 560898
rect 415794 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 416414 525454
rect 415794 525134 416414 525218
rect 415794 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 416414 525134
rect 415794 489454 416414 524898
rect 415794 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 416414 489454
rect 415794 489134 416414 489218
rect 415794 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 416414 489134
rect 415794 482000 416414 488898
rect 419514 673174 420134 707162
rect 419514 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 420134 673174
rect 419514 672854 420134 672938
rect 419514 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 420134 672854
rect 419514 637174 420134 672618
rect 419514 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 420134 637174
rect 419514 636854 420134 636938
rect 419514 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 420134 636854
rect 419514 601174 420134 636618
rect 419514 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 420134 601174
rect 419514 600854 420134 600938
rect 419514 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 420134 600854
rect 419514 565174 420134 600618
rect 419514 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 420134 565174
rect 419514 564854 420134 564938
rect 419514 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 420134 564854
rect 419514 529174 420134 564618
rect 419514 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 420134 529174
rect 419514 528854 420134 528938
rect 419514 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 420134 528854
rect 419514 493174 420134 528618
rect 419514 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 420134 493174
rect 419514 492854 420134 492938
rect 419514 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 420134 492854
rect 419514 482000 420134 492618
rect 423234 676894 423854 709082
rect 423234 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 423854 676894
rect 423234 676574 423854 676658
rect 423234 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 423854 676574
rect 423234 640894 423854 676338
rect 423234 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 423854 640894
rect 423234 640574 423854 640658
rect 423234 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 423854 640574
rect 423234 604894 423854 640338
rect 423234 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 423854 604894
rect 423234 604574 423854 604658
rect 423234 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 423854 604574
rect 423234 568894 423854 604338
rect 423234 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 423854 568894
rect 423234 568574 423854 568658
rect 423234 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 423854 568574
rect 423234 532894 423854 568338
rect 423234 532658 423266 532894
rect 423502 532658 423586 532894
rect 423822 532658 423854 532894
rect 423234 532574 423854 532658
rect 423234 532338 423266 532574
rect 423502 532338 423586 532574
rect 423822 532338 423854 532574
rect 423234 496894 423854 532338
rect 423234 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 423854 496894
rect 423234 496574 423854 496658
rect 423234 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 423854 496574
rect 423234 482000 423854 496338
rect 426954 680614 427574 711002
rect 444954 710598 445574 711590
rect 444954 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 445574 710598
rect 444954 710278 445574 710362
rect 444954 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 445574 710278
rect 441234 708678 441854 709670
rect 441234 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 441854 708678
rect 441234 708358 441854 708442
rect 441234 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 441854 708358
rect 437514 706758 438134 707750
rect 437514 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 438134 706758
rect 437514 706438 438134 706522
rect 437514 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 438134 706438
rect 426954 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 427574 680614
rect 426954 680294 427574 680378
rect 426954 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 427574 680294
rect 426954 644614 427574 680058
rect 426954 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 427574 644614
rect 426954 644294 427574 644378
rect 426954 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 427574 644294
rect 426954 608614 427574 644058
rect 426954 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 427574 608614
rect 426954 608294 427574 608378
rect 426954 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 427574 608294
rect 426954 572614 427574 608058
rect 426954 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 427574 572614
rect 426954 572294 427574 572378
rect 426954 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 427574 572294
rect 426954 536614 427574 572058
rect 426954 536378 426986 536614
rect 427222 536378 427306 536614
rect 427542 536378 427574 536614
rect 426954 536294 427574 536378
rect 426954 536058 426986 536294
rect 427222 536058 427306 536294
rect 427542 536058 427574 536294
rect 426954 500614 427574 536058
rect 426954 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 427574 500614
rect 426954 500294 427574 500378
rect 426954 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 427574 500294
rect 426954 482000 427574 500058
rect 433794 704838 434414 705830
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 482000 434414 506898
rect 437514 691174 438134 706202
rect 437514 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 438134 691174
rect 437514 690854 438134 690938
rect 437514 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 438134 690854
rect 437514 655174 438134 690618
rect 437514 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 438134 655174
rect 437514 654854 438134 654938
rect 437514 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 438134 654854
rect 437514 619174 438134 654618
rect 437514 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 438134 619174
rect 437514 618854 438134 618938
rect 437514 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 438134 618854
rect 437514 583174 438134 618618
rect 437514 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 438134 583174
rect 437514 582854 438134 582938
rect 437514 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 438134 582854
rect 437514 547174 438134 582618
rect 437514 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 438134 547174
rect 437514 546854 438134 546938
rect 437514 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 438134 546854
rect 437514 511174 438134 546618
rect 437514 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 438134 511174
rect 437514 510854 438134 510938
rect 437514 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 438134 510854
rect 437514 482000 438134 510618
rect 441234 694894 441854 708122
rect 441234 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 441854 694894
rect 441234 694574 441854 694658
rect 441234 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 441854 694574
rect 441234 658894 441854 694338
rect 441234 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 441854 658894
rect 441234 658574 441854 658658
rect 441234 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 441854 658574
rect 441234 622894 441854 658338
rect 441234 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 441854 622894
rect 441234 622574 441854 622658
rect 441234 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 441854 622574
rect 441234 586894 441854 622338
rect 441234 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 441854 586894
rect 441234 586574 441854 586658
rect 441234 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 441854 586574
rect 441234 550894 441854 586338
rect 441234 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 441854 550894
rect 441234 550574 441854 550658
rect 441234 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 441854 550574
rect 441234 514894 441854 550338
rect 441234 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 441854 514894
rect 441234 514574 441854 514658
rect 441234 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 441854 514574
rect 441234 482000 441854 514338
rect 444954 698614 445574 710042
rect 462954 711558 463574 711590
rect 462954 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 463574 711558
rect 462954 711238 463574 711322
rect 462954 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 463574 711238
rect 459234 709638 459854 709670
rect 459234 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 459854 709638
rect 459234 709318 459854 709402
rect 459234 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 459854 709318
rect 455514 707718 456134 707750
rect 455514 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 456134 707718
rect 455514 707398 456134 707482
rect 455514 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 456134 707398
rect 444954 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 445574 698614
rect 444954 698294 445574 698378
rect 444954 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 445574 698294
rect 444954 662614 445574 698058
rect 444954 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 445574 662614
rect 444954 662294 445574 662378
rect 444954 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 445574 662294
rect 444954 626614 445574 662058
rect 444954 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 445574 626614
rect 444954 626294 445574 626378
rect 444954 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 445574 626294
rect 444954 590614 445574 626058
rect 444954 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 445574 590614
rect 444954 590294 445574 590378
rect 444954 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 445574 590294
rect 444954 554614 445574 590058
rect 444954 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 445574 554614
rect 444954 554294 445574 554378
rect 444954 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 445574 554294
rect 444954 518614 445574 554058
rect 444954 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 445574 518614
rect 444954 518294 445574 518378
rect 444954 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 445574 518294
rect 444954 482614 445574 518058
rect 444954 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 445574 482614
rect 444954 482294 445574 482378
rect 444954 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 445574 482294
rect 444954 482000 445574 482058
rect 451794 705798 452414 705830
rect 451794 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 452414 705798
rect 451794 705478 452414 705562
rect 451794 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 452414 705478
rect 451794 669454 452414 705242
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 482000 452414 488898
rect 455514 673174 456134 707162
rect 455514 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 456134 673174
rect 455514 672854 456134 672938
rect 455514 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 456134 672854
rect 455514 637174 456134 672618
rect 455514 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 456134 637174
rect 455514 636854 456134 636938
rect 455514 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 456134 636854
rect 455514 601174 456134 636618
rect 455514 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 456134 601174
rect 455514 600854 456134 600938
rect 455514 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 456134 600854
rect 455514 565174 456134 600618
rect 455514 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 456134 565174
rect 455514 564854 456134 564938
rect 455514 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 456134 564854
rect 455514 529174 456134 564618
rect 455514 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 456134 529174
rect 455514 528854 456134 528938
rect 455514 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 456134 528854
rect 455514 493174 456134 528618
rect 455514 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 456134 493174
rect 455514 492854 456134 492938
rect 455514 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 456134 492854
rect 455514 482000 456134 492618
rect 459234 676894 459854 709082
rect 459234 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 459854 676894
rect 459234 676574 459854 676658
rect 459234 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 459854 676574
rect 459234 640894 459854 676338
rect 459234 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 459854 640894
rect 459234 640574 459854 640658
rect 459234 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 459854 640574
rect 459234 604894 459854 640338
rect 459234 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 459854 604894
rect 459234 604574 459854 604658
rect 459234 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 459854 604574
rect 459234 568894 459854 604338
rect 459234 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 459854 568894
rect 459234 568574 459854 568658
rect 459234 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 459854 568574
rect 459234 532894 459854 568338
rect 459234 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 459854 532894
rect 459234 532574 459854 532658
rect 459234 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 459854 532574
rect 459234 496894 459854 532338
rect 459234 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 459854 496894
rect 459234 496574 459854 496658
rect 459234 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 459854 496574
rect 459234 482000 459854 496338
rect 462954 680614 463574 711002
rect 480954 710598 481574 711590
rect 480954 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 481574 710598
rect 480954 710278 481574 710362
rect 480954 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 481574 710278
rect 477234 708678 477854 709670
rect 477234 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 477854 708678
rect 477234 708358 477854 708442
rect 477234 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 477854 708358
rect 473514 706758 474134 707750
rect 473514 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 474134 706758
rect 473514 706438 474134 706522
rect 473514 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 474134 706438
rect 462954 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 463574 680614
rect 462954 680294 463574 680378
rect 462954 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 463574 680294
rect 462954 644614 463574 680058
rect 462954 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 463574 644614
rect 462954 644294 463574 644378
rect 462954 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 463574 644294
rect 462954 608614 463574 644058
rect 462954 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 463574 608614
rect 462954 608294 463574 608378
rect 462954 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 463574 608294
rect 462954 572614 463574 608058
rect 462954 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 463574 572614
rect 462954 572294 463574 572378
rect 462954 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 463574 572294
rect 462954 536614 463574 572058
rect 462954 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 463574 536614
rect 462954 536294 463574 536378
rect 462954 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 463574 536294
rect 462954 500614 463574 536058
rect 462954 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 463574 500614
rect 462954 500294 463574 500378
rect 462954 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 463574 500294
rect 462954 482000 463574 500058
rect 469794 704838 470414 705830
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 482000 470414 506898
rect 473514 691174 474134 706202
rect 473514 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 474134 691174
rect 473514 690854 474134 690938
rect 473514 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 474134 690854
rect 473514 655174 474134 690618
rect 473514 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 474134 655174
rect 473514 654854 474134 654938
rect 473514 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 474134 654854
rect 473514 619174 474134 654618
rect 473514 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 474134 619174
rect 473514 618854 474134 618938
rect 473514 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 474134 618854
rect 473514 583174 474134 618618
rect 473514 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 474134 583174
rect 473514 582854 474134 582938
rect 473514 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 474134 582854
rect 473514 547174 474134 582618
rect 473514 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 474134 547174
rect 473514 546854 474134 546938
rect 473514 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 474134 546854
rect 473514 511174 474134 546618
rect 473514 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 474134 511174
rect 473514 510854 474134 510938
rect 473514 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 474134 510854
rect 473514 482000 474134 510618
rect 477234 694894 477854 708122
rect 477234 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 477854 694894
rect 477234 694574 477854 694658
rect 477234 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 477854 694574
rect 477234 658894 477854 694338
rect 477234 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 477854 658894
rect 477234 658574 477854 658658
rect 477234 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 477854 658574
rect 477234 622894 477854 658338
rect 477234 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 477854 622894
rect 477234 622574 477854 622658
rect 477234 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 477854 622574
rect 477234 586894 477854 622338
rect 477234 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 477854 586894
rect 477234 586574 477854 586658
rect 477234 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 477854 586574
rect 477234 550894 477854 586338
rect 477234 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 477854 550894
rect 477234 550574 477854 550658
rect 477234 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 477854 550574
rect 477234 514894 477854 550338
rect 477234 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 477854 514894
rect 477234 514574 477854 514658
rect 477234 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 477854 514574
rect 477234 482000 477854 514338
rect 480954 698614 481574 710042
rect 498954 711558 499574 711590
rect 498954 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 499574 711558
rect 498954 711238 499574 711322
rect 498954 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 499574 711238
rect 495234 709638 495854 709670
rect 495234 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 495854 709638
rect 495234 709318 495854 709402
rect 495234 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 495854 709318
rect 491514 707718 492134 707750
rect 491514 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 492134 707718
rect 491514 707398 492134 707482
rect 491514 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 492134 707398
rect 480954 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 481574 698614
rect 480954 698294 481574 698378
rect 480954 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 481574 698294
rect 480954 662614 481574 698058
rect 480954 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 481574 662614
rect 480954 662294 481574 662378
rect 480954 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 481574 662294
rect 480954 626614 481574 662058
rect 480954 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 481574 626614
rect 480954 626294 481574 626378
rect 480954 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 481574 626294
rect 480954 590614 481574 626058
rect 480954 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 481574 590614
rect 480954 590294 481574 590378
rect 480954 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 481574 590294
rect 480954 554614 481574 590058
rect 480954 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 481574 554614
rect 480954 554294 481574 554378
rect 480954 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 481574 554294
rect 480954 518614 481574 554058
rect 480954 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 481574 518614
rect 480954 518294 481574 518378
rect 480954 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 481574 518294
rect 480954 482614 481574 518058
rect 480954 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 481574 482614
rect 480954 482294 481574 482378
rect 480954 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 481574 482294
rect 480954 482000 481574 482058
rect 487794 705798 488414 705830
rect 487794 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 488414 705798
rect 487794 705478 488414 705562
rect 487794 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 488414 705478
rect 487794 669454 488414 705242
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 561454 488414 596898
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 482000 488414 488898
rect 491514 673174 492134 707162
rect 491514 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 492134 673174
rect 491514 672854 492134 672938
rect 491514 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 492134 672854
rect 491514 637174 492134 672618
rect 491514 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 492134 637174
rect 491514 636854 492134 636938
rect 491514 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 492134 636854
rect 491514 601174 492134 636618
rect 491514 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 492134 601174
rect 491514 600854 492134 600938
rect 491514 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 492134 600854
rect 491514 565174 492134 600618
rect 491514 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 492134 565174
rect 491514 564854 492134 564938
rect 491514 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 492134 564854
rect 491514 529174 492134 564618
rect 491514 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 492134 529174
rect 491514 528854 492134 528938
rect 491514 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 492134 528854
rect 491514 493174 492134 528618
rect 491514 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 492134 493174
rect 491514 492854 492134 492938
rect 491514 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 492134 492854
rect 491514 482000 492134 492618
rect 495234 676894 495854 709082
rect 495234 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 495854 676894
rect 495234 676574 495854 676658
rect 495234 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 495854 676574
rect 495234 640894 495854 676338
rect 495234 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 495854 640894
rect 495234 640574 495854 640658
rect 495234 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 495854 640574
rect 495234 604894 495854 640338
rect 495234 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 495854 604894
rect 495234 604574 495854 604658
rect 495234 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 495854 604574
rect 495234 568894 495854 604338
rect 495234 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 495854 568894
rect 495234 568574 495854 568658
rect 495234 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 495854 568574
rect 495234 532894 495854 568338
rect 495234 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 495854 532894
rect 495234 532574 495854 532658
rect 495234 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 495854 532574
rect 495234 496894 495854 532338
rect 495234 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 495854 496894
rect 495234 496574 495854 496658
rect 495234 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 495854 496574
rect 495234 482000 495854 496338
rect 498954 680614 499574 711002
rect 516954 710598 517574 711590
rect 516954 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 517574 710598
rect 516954 710278 517574 710362
rect 516954 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 517574 710278
rect 513234 708678 513854 709670
rect 513234 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 513854 708678
rect 513234 708358 513854 708442
rect 513234 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 513854 708358
rect 509514 706758 510134 707750
rect 509514 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 510134 706758
rect 509514 706438 510134 706522
rect 509514 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 510134 706438
rect 498954 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 499574 680614
rect 498954 680294 499574 680378
rect 498954 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 499574 680294
rect 498954 644614 499574 680058
rect 498954 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 499574 644614
rect 498954 644294 499574 644378
rect 498954 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 499574 644294
rect 498954 608614 499574 644058
rect 498954 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 499574 608614
rect 498954 608294 499574 608378
rect 498954 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 499574 608294
rect 498954 572614 499574 608058
rect 498954 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 499574 572614
rect 498954 572294 499574 572378
rect 498954 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 499574 572294
rect 498954 536614 499574 572058
rect 498954 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 499574 536614
rect 498954 536294 499574 536378
rect 498954 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 499574 536294
rect 498954 500614 499574 536058
rect 498954 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 499574 500614
rect 498954 500294 499574 500378
rect 498954 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 499574 500294
rect 498954 482000 499574 500058
rect 505794 704838 506414 705830
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 482000 506414 506898
rect 509514 691174 510134 706202
rect 509514 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 510134 691174
rect 509514 690854 510134 690938
rect 509514 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 510134 690854
rect 509514 655174 510134 690618
rect 509514 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 510134 655174
rect 509514 654854 510134 654938
rect 509514 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 510134 654854
rect 509514 619174 510134 654618
rect 509514 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 510134 619174
rect 509514 618854 510134 618938
rect 509514 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 510134 618854
rect 509514 583174 510134 618618
rect 509514 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 510134 583174
rect 509514 582854 510134 582938
rect 509514 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 510134 582854
rect 509514 547174 510134 582618
rect 509514 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 510134 547174
rect 509514 546854 510134 546938
rect 509514 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 510134 546854
rect 509514 511174 510134 546618
rect 509514 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 510134 511174
rect 509514 510854 510134 510938
rect 509514 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 510134 510854
rect 509514 482000 510134 510618
rect 513234 694894 513854 708122
rect 513234 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 513854 694894
rect 513234 694574 513854 694658
rect 513234 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 513854 694574
rect 513234 658894 513854 694338
rect 513234 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 513854 658894
rect 513234 658574 513854 658658
rect 513234 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 513854 658574
rect 513234 622894 513854 658338
rect 513234 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 513854 622894
rect 513234 622574 513854 622658
rect 513234 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 513854 622574
rect 513234 586894 513854 622338
rect 513234 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 513854 586894
rect 513234 586574 513854 586658
rect 513234 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 513854 586574
rect 513234 550894 513854 586338
rect 513234 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 513854 550894
rect 513234 550574 513854 550658
rect 513234 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 513854 550574
rect 513234 514894 513854 550338
rect 513234 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 513854 514894
rect 513234 514574 513854 514658
rect 513234 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 513854 514574
rect 513234 482000 513854 514338
rect 516954 698614 517574 710042
rect 534954 711558 535574 711590
rect 534954 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 535574 711558
rect 534954 711238 535574 711322
rect 534954 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 535574 711238
rect 531234 709638 531854 709670
rect 531234 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 531854 709638
rect 531234 709318 531854 709402
rect 531234 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 531854 709318
rect 527514 707718 528134 707750
rect 527514 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 528134 707718
rect 527514 707398 528134 707482
rect 527514 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 528134 707398
rect 516954 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 517574 698614
rect 516954 698294 517574 698378
rect 516954 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 517574 698294
rect 516954 662614 517574 698058
rect 516954 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 517574 662614
rect 516954 662294 517574 662378
rect 516954 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 517574 662294
rect 516954 626614 517574 662058
rect 516954 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 517574 626614
rect 516954 626294 517574 626378
rect 516954 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 517574 626294
rect 516954 590614 517574 626058
rect 516954 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 517574 590614
rect 516954 590294 517574 590378
rect 516954 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 517574 590294
rect 516954 554614 517574 590058
rect 516954 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 517574 554614
rect 516954 554294 517574 554378
rect 516954 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 517574 554294
rect 516954 518614 517574 554058
rect 516954 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 517574 518614
rect 516954 518294 517574 518378
rect 516954 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 517574 518294
rect 516954 482614 517574 518058
rect 516954 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 517574 482614
rect 516954 482294 517574 482378
rect 516954 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 517574 482294
rect 516954 482000 517574 482058
rect 523794 705798 524414 705830
rect 523794 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 524414 705798
rect 523794 705478 524414 705562
rect 523794 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 524414 705478
rect 523794 669454 524414 705242
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 482000 524414 488898
rect 527514 673174 528134 707162
rect 527514 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 528134 673174
rect 527514 672854 528134 672938
rect 527514 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 528134 672854
rect 527514 637174 528134 672618
rect 527514 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 528134 637174
rect 527514 636854 528134 636938
rect 527514 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 528134 636854
rect 527514 601174 528134 636618
rect 527514 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 528134 601174
rect 527514 600854 528134 600938
rect 527514 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 528134 600854
rect 527514 565174 528134 600618
rect 527514 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 528134 565174
rect 527514 564854 528134 564938
rect 527514 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 528134 564854
rect 527514 529174 528134 564618
rect 527514 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 528134 529174
rect 527514 528854 528134 528938
rect 527514 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 528134 528854
rect 527514 493174 528134 528618
rect 527514 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 528134 493174
rect 527514 492854 528134 492938
rect 527514 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 528134 492854
rect 527514 482000 528134 492618
rect 531234 676894 531854 709082
rect 531234 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 531854 676894
rect 531234 676574 531854 676658
rect 531234 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 531854 676574
rect 531234 640894 531854 676338
rect 531234 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 531854 640894
rect 531234 640574 531854 640658
rect 531234 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 531854 640574
rect 531234 604894 531854 640338
rect 531234 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 531854 604894
rect 531234 604574 531854 604658
rect 531234 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 531854 604574
rect 531234 568894 531854 604338
rect 531234 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 531854 568894
rect 531234 568574 531854 568658
rect 531234 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 531854 568574
rect 531234 532894 531854 568338
rect 531234 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 531854 532894
rect 531234 532574 531854 532658
rect 531234 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 531854 532574
rect 531234 496894 531854 532338
rect 531234 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 531854 496894
rect 531234 496574 531854 496658
rect 531234 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 531854 496574
rect 531234 482000 531854 496338
rect 534954 680614 535574 711002
rect 552954 710598 553574 711590
rect 552954 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 553574 710598
rect 552954 710278 553574 710362
rect 552954 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 553574 710278
rect 549234 708678 549854 709670
rect 549234 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 549854 708678
rect 549234 708358 549854 708442
rect 549234 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 549854 708358
rect 545514 706758 546134 707750
rect 545514 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 546134 706758
rect 545514 706438 546134 706522
rect 545514 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 546134 706438
rect 534954 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 535574 680614
rect 534954 680294 535574 680378
rect 534954 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 535574 680294
rect 534954 644614 535574 680058
rect 534954 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 535574 644614
rect 534954 644294 535574 644378
rect 534954 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 535574 644294
rect 534954 608614 535574 644058
rect 534954 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 535574 608614
rect 534954 608294 535574 608378
rect 534954 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 535574 608294
rect 534954 572614 535574 608058
rect 541794 704838 542414 705830
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 536787 596868 536853 596869
rect 536787 596804 536788 596868
rect 536852 596804 536853 596868
rect 536787 596803 536853 596804
rect 534954 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 535574 572614
rect 534954 572294 535574 572378
rect 534954 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 535574 572294
rect 534954 536614 535574 572058
rect 534954 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 535574 536614
rect 534954 536294 535574 536378
rect 534954 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 535574 536294
rect 534954 500614 535574 536058
rect 534954 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 535574 500614
rect 534954 500294 535574 500378
rect 534954 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 535574 500294
rect 534954 482000 535574 500058
rect 244208 471454 244528 471486
rect 244208 471218 244250 471454
rect 244486 471218 244528 471454
rect 244208 471134 244528 471218
rect 244208 470898 244250 471134
rect 244486 470898 244528 471134
rect 244208 470866 244528 470898
rect 274928 471454 275248 471486
rect 274928 471218 274970 471454
rect 275206 471218 275248 471454
rect 274928 471134 275248 471218
rect 274928 470898 274970 471134
rect 275206 470898 275248 471134
rect 274928 470866 275248 470898
rect 305648 471454 305968 471486
rect 305648 471218 305690 471454
rect 305926 471218 305968 471454
rect 305648 471134 305968 471218
rect 305648 470898 305690 471134
rect 305926 470898 305968 471134
rect 305648 470866 305968 470898
rect 336368 471454 336688 471486
rect 336368 471218 336410 471454
rect 336646 471218 336688 471454
rect 336368 471134 336688 471218
rect 336368 470898 336410 471134
rect 336646 470898 336688 471134
rect 336368 470866 336688 470898
rect 367088 471454 367408 471486
rect 367088 471218 367130 471454
rect 367366 471218 367408 471454
rect 367088 471134 367408 471218
rect 367088 470898 367130 471134
rect 367366 470898 367408 471134
rect 367088 470866 367408 470898
rect 397808 471454 398128 471486
rect 397808 471218 397850 471454
rect 398086 471218 398128 471454
rect 397808 471134 398128 471218
rect 397808 470898 397850 471134
rect 398086 470898 398128 471134
rect 397808 470866 398128 470898
rect 428528 471454 428848 471486
rect 428528 471218 428570 471454
rect 428806 471218 428848 471454
rect 428528 471134 428848 471218
rect 428528 470898 428570 471134
rect 428806 470898 428848 471134
rect 428528 470866 428848 470898
rect 459248 471454 459568 471486
rect 459248 471218 459290 471454
rect 459526 471218 459568 471454
rect 459248 471134 459568 471218
rect 459248 470898 459290 471134
rect 459526 470898 459568 471134
rect 459248 470866 459568 470898
rect 489968 471454 490288 471486
rect 489968 471218 490010 471454
rect 490246 471218 490288 471454
rect 489968 471134 490288 471218
rect 489968 470898 490010 471134
rect 490246 470898 490288 471134
rect 489968 470866 490288 470898
rect 520688 471454 521008 471486
rect 520688 471218 520730 471454
rect 520966 471218 521008 471454
rect 520688 471134 521008 471218
rect 520688 470898 520730 471134
rect 520966 470898 521008 471134
rect 520688 470866 521008 470898
rect 259568 453454 259888 453486
rect 259568 453218 259610 453454
rect 259846 453218 259888 453454
rect 259568 453134 259888 453218
rect 259568 452898 259610 453134
rect 259846 452898 259888 453134
rect 259568 452866 259888 452898
rect 290288 453454 290608 453486
rect 290288 453218 290330 453454
rect 290566 453218 290608 453454
rect 290288 453134 290608 453218
rect 290288 452898 290330 453134
rect 290566 452898 290608 453134
rect 290288 452866 290608 452898
rect 321008 453454 321328 453486
rect 321008 453218 321050 453454
rect 321286 453218 321328 453454
rect 321008 453134 321328 453218
rect 321008 452898 321050 453134
rect 321286 452898 321328 453134
rect 321008 452866 321328 452898
rect 351728 453454 352048 453486
rect 351728 453218 351770 453454
rect 352006 453218 352048 453454
rect 351728 453134 352048 453218
rect 351728 452898 351770 453134
rect 352006 452898 352048 453134
rect 351728 452866 352048 452898
rect 382448 453454 382768 453486
rect 382448 453218 382490 453454
rect 382726 453218 382768 453454
rect 382448 453134 382768 453218
rect 382448 452898 382490 453134
rect 382726 452898 382768 453134
rect 382448 452866 382768 452898
rect 413168 453454 413488 453486
rect 413168 453218 413210 453454
rect 413446 453218 413488 453454
rect 413168 453134 413488 453218
rect 413168 452898 413210 453134
rect 413446 452898 413488 453134
rect 413168 452866 413488 452898
rect 443888 453454 444208 453486
rect 443888 453218 443930 453454
rect 444166 453218 444208 453454
rect 443888 453134 444208 453218
rect 443888 452898 443930 453134
rect 444166 452898 444208 453134
rect 443888 452866 444208 452898
rect 474608 453454 474928 453486
rect 474608 453218 474650 453454
rect 474886 453218 474928 453454
rect 474608 453134 474928 453218
rect 474608 452898 474650 453134
rect 474886 452898 474928 453134
rect 474608 452866 474928 452898
rect 505328 453454 505648 453486
rect 505328 453218 505370 453454
rect 505606 453218 505648 453454
rect 505328 453134 505648 453218
rect 505328 452898 505370 453134
rect 505606 452898 505648 453134
rect 505328 452866 505648 452898
rect 536048 453454 536368 453486
rect 536048 453218 536090 453454
rect 536326 453218 536368 453454
rect 536048 453134 536368 453218
rect 536048 452898 536090 453134
rect 536326 452898 536368 453134
rect 536048 452866 536368 452898
rect 244208 435454 244528 435486
rect 244208 435218 244250 435454
rect 244486 435218 244528 435454
rect 244208 435134 244528 435218
rect 244208 434898 244250 435134
rect 244486 434898 244528 435134
rect 244208 434866 244528 434898
rect 274928 435454 275248 435486
rect 274928 435218 274970 435454
rect 275206 435218 275248 435454
rect 274928 435134 275248 435218
rect 274928 434898 274970 435134
rect 275206 434898 275248 435134
rect 274928 434866 275248 434898
rect 305648 435454 305968 435486
rect 305648 435218 305690 435454
rect 305926 435218 305968 435454
rect 305648 435134 305968 435218
rect 305648 434898 305690 435134
rect 305926 434898 305968 435134
rect 305648 434866 305968 434898
rect 336368 435454 336688 435486
rect 336368 435218 336410 435454
rect 336646 435218 336688 435454
rect 336368 435134 336688 435218
rect 336368 434898 336410 435134
rect 336646 434898 336688 435134
rect 336368 434866 336688 434898
rect 367088 435454 367408 435486
rect 367088 435218 367130 435454
rect 367366 435218 367408 435454
rect 367088 435134 367408 435218
rect 367088 434898 367130 435134
rect 367366 434898 367408 435134
rect 367088 434866 367408 434898
rect 397808 435454 398128 435486
rect 397808 435218 397850 435454
rect 398086 435218 398128 435454
rect 397808 435134 398128 435218
rect 397808 434898 397850 435134
rect 398086 434898 398128 435134
rect 397808 434866 398128 434898
rect 428528 435454 428848 435486
rect 428528 435218 428570 435454
rect 428806 435218 428848 435454
rect 428528 435134 428848 435218
rect 428528 434898 428570 435134
rect 428806 434898 428848 435134
rect 428528 434866 428848 434898
rect 459248 435454 459568 435486
rect 459248 435218 459290 435454
rect 459526 435218 459568 435454
rect 459248 435134 459568 435218
rect 459248 434898 459290 435134
rect 459526 434898 459568 435134
rect 459248 434866 459568 434898
rect 489968 435454 490288 435486
rect 489968 435218 490010 435454
rect 490246 435218 490288 435454
rect 489968 435134 490288 435218
rect 489968 434898 490010 435134
rect 490246 434898 490288 435134
rect 489968 434866 490288 434898
rect 520688 435454 521008 435486
rect 520688 435218 520730 435454
rect 520966 435218 521008 435454
rect 520688 435134 521008 435218
rect 520688 434898 520730 435134
rect 520966 434898 521008 435134
rect 520688 434866 521008 434898
rect 259568 417454 259888 417486
rect 259568 417218 259610 417454
rect 259846 417218 259888 417454
rect 259568 417134 259888 417218
rect 259568 416898 259610 417134
rect 259846 416898 259888 417134
rect 259568 416866 259888 416898
rect 290288 417454 290608 417486
rect 290288 417218 290330 417454
rect 290566 417218 290608 417454
rect 290288 417134 290608 417218
rect 290288 416898 290330 417134
rect 290566 416898 290608 417134
rect 290288 416866 290608 416898
rect 321008 417454 321328 417486
rect 321008 417218 321050 417454
rect 321286 417218 321328 417454
rect 321008 417134 321328 417218
rect 321008 416898 321050 417134
rect 321286 416898 321328 417134
rect 321008 416866 321328 416898
rect 351728 417454 352048 417486
rect 351728 417218 351770 417454
rect 352006 417218 352048 417454
rect 351728 417134 352048 417218
rect 351728 416898 351770 417134
rect 352006 416898 352048 417134
rect 351728 416866 352048 416898
rect 382448 417454 382768 417486
rect 382448 417218 382490 417454
rect 382726 417218 382768 417454
rect 382448 417134 382768 417218
rect 382448 416898 382490 417134
rect 382726 416898 382768 417134
rect 382448 416866 382768 416898
rect 413168 417454 413488 417486
rect 413168 417218 413210 417454
rect 413446 417218 413488 417454
rect 413168 417134 413488 417218
rect 413168 416898 413210 417134
rect 413446 416898 413488 417134
rect 413168 416866 413488 416898
rect 443888 417454 444208 417486
rect 443888 417218 443930 417454
rect 444166 417218 444208 417454
rect 443888 417134 444208 417218
rect 443888 416898 443930 417134
rect 444166 416898 444208 417134
rect 443888 416866 444208 416898
rect 474608 417454 474928 417486
rect 474608 417218 474650 417454
rect 474886 417218 474928 417454
rect 474608 417134 474928 417218
rect 474608 416898 474650 417134
rect 474886 416898 474928 417134
rect 474608 416866 474928 416898
rect 505328 417454 505648 417486
rect 505328 417218 505370 417454
rect 505606 417218 505648 417454
rect 505328 417134 505648 417218
rect 505328 416898 505370 417134
rect 505606 416898 505648 417134
rect 505328 416866 505648 416898
rect 536048 417454 536368 417486
rect 536048 417218 536090 417454
rect 536326 417218 536368 417454
rect 536048 417134 536368 417218
rect 536048 416898 536090 417134
rect 536326 416898 536368 417134
rect 536048 416866 536368 416898
rect 244208 399454 244528 399486
rect 244208 399218 244250 399454
rect 244486 399218 244528 399454
rect 244208 399134 244528 399218
rect 244208 398898 244250 399134
rect 244486 398898 244528 399134
rect 244208 398866 244528 398898
rect 274928 399454 275248 399486
rect 274928 399218 274970 399454
rect 275206 399218 275248 399454
rect 274928 399134 275248 399218
rect 274928 398898 274970 399134
rect 275206 398898 275248 399134
rect 274928 398866 275248 398898
rect 305648 399454 305968 399486
rect 305648 399218 305690 399454
rect 305926 399218 305968 399454
rect 305648 399134 305968 399218
rect 305648 398898 305690 399134
rect 305926 398898 305968 399134
rect 305648 398866 305968 398898
rect 336368 399454 336688 399486
rect 336368 399218 336410 399454
rect 336646 399218 336688 399454
rect 336368 399134 336688 399218
rect 336368 398898 336410 399134
rect 336646 398898 336688 399134
rect 336368 398866 336688 398898
rect 367088 399454 367408 399486
rect 367088 399218 367130 399454
rect 367366 399218 367408 399454
rect 367088 399134 367408 399218
rect 367088 398898 367130 399134
rect 367366 398898 367408 399134
rect 367088 398866 367408 398898
rect 397808 399454 398128 399486
rect 397808 399218 397850 399454
rect 398086 399218 398128 399454
rect 397808 399134 398128 399218
rect 397808 398898 397850 399134
rect 398086 398898 398128 399134
rect 397808 398866 398128 398898
rect 428528 399454 428848 399486
rect 428528 399218 428570 399454
rect 428806 399218 428848 399454
rect 428528 399134 428848 399218
rect 428528 398898 428570 399134
rect 428806 398898 428848 399134
rect 428528 398866 428848 398898
rect 459248 399454 459568 399486
rect 459248 399218 459290 399454
rect 459526 399218 459568 399454
rect 459248 399134 459568 399218
rect 459248 398898 459290 399134
rect 459526 398898 459568 399134
rect 459248 398866 459568 398898
rect 489968 399454 490288 399486
rect 489968 399218 490010 399454
rect 490246 399218 490288 399454
rect 489968 399134 490288 399218
rect 489968 398898 490010 399134
rect 490246 398898 490288 399134
rect 489968 398866 490288 398898
rect 520688 399454 521008 399486
rect 520688 399218 520730 399454
rect 520966 399218 521008 399454
rect 520688 399134 521008 399218
rect 520688 398898 520730 399134
rect 520966 398898 521008 399134
rect 520688 398866 521008 398898
rect 259568 381454 259888 381486
rect 259568 381218 259610 381454
rect 259846 381218 259888 381454
rect 259568 381134 259888 381218
rect 259568 380898 259610 381134
rect 259846 380898 259888 381134
rect 259568 380866 259888 380898
rect 290288 381454 290608 381486
rect 290288 381218 290330 381454
rect 290566 381218 290608 381454
rect 290288 381134 290608 381218
rect 290288 380898 290330 381134
rect 290566 380898 290608 381134
rect 290288 380866 290608 380898
rect 321008 381454 321328 381486
rect 321008 381218 321050 381454
rect 321286 381218 321328 381454
rect 321008 381134 321328 381218
rect 321008 380898 321050 381134
rect 321286 380898 321328 381134
rect 321008 380866 321328 380898
rect 351728 381454 352048 381486
rect 351728 381218 351770 381454
rect 352006 381218 352048 381454
rect 351728 381134 352048 381218
rect 351728 380898 351770 381134
rect 352006 380898 352048 381134
rect 351728 380866 352048 380898
rect 382448 381454 382768 381486
rect 382448 381218 382490 381454
rect 382726 381218 382768 381454
rect 382448 381134 382768 381218
rect 382448 380898 382490 381134
rect 382726 380898 382768 381134
rect 382448 380866 382768 380898
rect 413168 381454 413488 381486
rect 413168 381218 413210 381454
rect 413446 381218 413488 381454
rect 413168 381134 413488 381218
rect 413168 380898 413210 381134
rect 413446 380898 413488 381134
rect 413168 380866 413488 380898
rect 443888 381454 444208 381486
rect 443888 381218 443930 381454
rect 444166 381218 444208 381454
rect 443888 381134 444208 381218
rect 443888 380898 443930 381134
rect 444166 380898 444208 381134
rect 443888 380866 444208 380898
rect 474608 381454 474928 381486
rect 474608 381218 474650 381454
rect 474886 381218 474928 381454
rect 474608 381134 474928 381218
rect 474608 380898 474650 381134
rect 474886 380898 474928 381134
rect 474608 380866 474928 380898
rect 505328 381454 505648 381486
rect 505328 381218 505370 381454
rect 505606 381218 505648 381454
rect 505328 381134 505648 381218
rect 505328 380898 505370 381134
rect 505606 380898 505648 381134
rect 505328 380866 505648 380898
rect 536048 381454 536368 381486
rect 536048 381218 536090 381454
rect 536326 381218 536368 381454
rect 536048 381134 536368 381218
rect 536048 380898 536090 381134
rect 536326 380898 536368 381134
rect 536048 380866 536368 380898
rect 244208 363454 244528 363486
rect 244208 363218 244250 363454
rect 244486 363218 244528 363454
rect 244208 363134 244528 363218
rect 244208 362898 244250 363134
rect 244486 362898 244528 363134
rect 244208 362866 244528 362898
rect 274928 363454 275248 363486
rect 274928 363218 274970 363454
rect 275206 363218 275248 363454
rect 274928 363134 275248 363218
rect 274928 362898 274970 363134
rect 275206 362898 275248 363134
rect 274928 362866 275248 362898
rect 305648 363454 305968 363486
rect 305648 363218 305690 363454
rect 305926 363218 305968 363454
rect 305648 363134 305968 363218
rect 305648 362898 305690 363134
rect 305926 362898 305968 363134
rect 305648 362866 305968 362898
rect 336368 363454 336688 363486
rect 336368 363218 336410 363454
rect 336646 363218 336688 363454
rect 336368 363134 336688 363218
rect 336368 362898 336410 363134
rect 336646 362898 336688 363134
rect 336368 362866 336688 362898
rect 367088 363454 367408 363486
rect 367088 363218 367130 363454
rect 367366 363218 367408 363454
rect 367088 363134 367408 363218
rect 367088 362898 367130 363134
rect 367366 362898 367408 363134
rect 367088 362866 367408 362898
rect 397808 363454 398128 363486
rect 397808 363218 397850 363454
rect 398086 363218 398128 363454
rect 397808 363134 398128 363218
rect 397808 362898 397850 363134
rect 398086 362898 398128 363134
rect 397808 362866 398128 362898
rect 428528 363454 428848 363486
rect 428528 363218 428570 363454
rect 428806 363218 428848 363454
rect 428528 363134 428848 363218
rect 428528 362898 428570 363134
rect 428806 362898 428848 363134
rect 428528 362866 428848 362898
rect 459248 363454 459568 363486
rect 459248 363218 459290 363454
rect 459526 363218 459568 363454
rect 459248 363134 459568 363218
rect 459248 362898 459290 363134
rect 459526 362898 459568 363134
rect 459248 362866 459568 362898
rect 489968 363454 490288 363486
rect 489968 363218 490010 363454
rect 490246 363218 490288 363454
rect 489968 363134 490288 363218
rect 489968 362898 490010 363134
rect 490246 362898 490288 363134
rect 489968 362866 490288 362898
rect 520688 363454 521008 363486
rect 520688 363218 520730 363454
rect 520966 363218 521008 363454
rect 520688 363134 521008 363218
rect 520688 362898 520730 363134
rect 520966 362898 521008 363134
rect 520688 362866 521008 362898
rect 259568 345454 259888 345486
rect 259568 345218 259610 345454
rect 259846 345218 259888 345454
rect 259568 345134 259888 345218
rect 259568 344898 259610 345134
rect 259846 344898 259888 345134
rect 259568 344866 259888 344898
rect 290288 345454 290608 345486
rect 290288 345218 290330 345454
rect 290566 345218 290608 345454
rect 290288 345134 290608 345218
rect 290288 344898 290330 345134
rect 290566 344898 290608 345134
rect 290288 344866 290608 344898
rect 321008 345454 321328 345486
rect 321008 345218 321050 345454
rect 321286 345218 321328 345454
rect 321008 345134 321328 345218
rect 321008 344898 321050 345134
rect 321286 344898 321328 345134
rect 321008 344866 321328 344898
rect 351728 345454 352048 345486
rect 351728 345218 351770 345454
rect 352006 345218 352048 345454
rect 351728 345134 352048 345218
rect 351728 344898 351770 345134
rect 352006 344898 352048 345134
rect 351728 344866 352048 344898
rect 382448 345454 382768 345486
rect 382448 345218 382490 345454
rect 382726 345218 382768 345454
rect 382448 345134 382768 345218
rect 382448 344898 382490 345134
rect 382726 344898 382768 345134
rect 382448 344866 382768 344898
rect 413168 345454 413488 345486
rect 413168 345218 413210 345454
rect 413446 345218 413488 345454
rect 413168 345134 413488 345218
rect 413168 344898 413210 345134
rect 413446 344898 413488 345134
rect 413168 344866 413488 344898
rect 443888 345454 444208 345486
rect 443888 345218 443930 345454
rect 444166 345218 444208 345454
rect 443888 345134 444208 345218
rect 443888 344898 443930 345134
rect 444166 344898 444208 345134
rect 443888 344866 444208 344898
rect 474608 345454 474928 345486
rect 474608 345218 474650 345454
rect 474886 345218 474928 345454
rect 474608 345134 474928 345218
rect 474608 344898 474650 345134
rect 474886 344898 474928 345134
rect 474608 344866 474928 344898
rect 505328 345454 505648 345486
rect 505328 345218 505370 345454
rect 505606 345218 505648 345454
rect 505328 345134 505648 345218
rect 505328 344898 505370 345134
rect 505606 344898 505648 345134
rect 505328 344866 505648 344898
rect 536048 345454 536368 345486
rect 536048 345218 536090 345454
rect 536326 345218 536368 345454
rect 536048 345134 536368 345218
rect 536048 344898 536090 345134
rect 536326 344898 536368 345134
rect 536048 344866 536368 344898
rect 244208 327454 244528 327486
rect 244208 327218 244250 327454
rect 244486 327218 244528 327454
rect 244208 327134 244528 327218
rect 244208 326898 244250 327134
rect 244486 326898 244528 327134
rect 244208 326866 244528 326898
rect 274928 327454 275248 327486
rect 274928 327218 274970 327454
rect 275206 327218 275248 327454
rect 274928 327134 275248 327218
rect 274928 326898 274970 327134
rect 275206 326898 275248 327134
rect 274928 326866 275248 326898
rect 305648 327454 305968 327486
rect 305648 327218 305690 327454
rect 305926 327218 305968 327454
rect 305648 327134 305968 327218
rect 305648 326898 305690 327134
rect 305926 326898 305968 327134
rect 305648 326866 305968 326898
rect 336368 327454 336688 327486
rect 336368 327218 336410 327454
rect 336646 327218 336688 327454
rect 336368 327134 336688 327218
rect 336368 326898 336410 327134
rect 336646 326898 336688 327134
rect 336368 326866 336688 326898
rect 367088 327454 367408 327486
rect 367088 327218 367130 327454
rect 367366 327218 367408 327454
rect 367088 327134 367408 327218
rect 367088 326898 367130 327134
rect 367366 326898 367408 327134
rect 367088 326866 367408 326898
rect 397808 327454 398128 327486
rect 397808 327218 397850 327454
rect 398086 327218 398128 327454
rect 397808 327134 398128 327218
rect 397808 326898 397850 327134
rect 398086 326898 398128 327134
rect 397808 326866 398128 326898
rect 428528 327454 428848 327486
rect 428528 327218 428570 327454
rect 428806 327218 428848 327454
rect 428528 327134 428848 327218
rect 428528 326898 428570 327134
rect 428806 326898 428848 327134
rect 428528 326866 428848 326898
rect 459248 327454 459568 327486
rect 459248 327218 459290 327454
rect 459526 327218 459568 327454
rect 459248 327134 459568 327218
rect 459248 326898 459290 327134
rect 459526 326898 459568 327134
rect 459248 326866 459568 326898
rect 489968 327454 490288 327486
rect 489968 327218 490010 327454
rect 490246 327218 490288 327454
rect 489968 327134 490288 327218
rect 489968 326898 490010 327134
rect 490246 326898 490288 327134
rect 489968 326866 490288 326898
rect 520688 327454 521008 327486
rect 520688 327218 520730 327454
rect 520966 327218 521008 327454
rect 520688 327134 521008 327218
rect 520688 326898 520730 327134
rect 520966 326898 521008 327134
rect 520688 326866 521008 326898
rect 259568 309454 259888 309486
rect 259568 309218 259610 309454
rect 259846 309218 259888 309454
rect 259568 309134 259888 309218
rect 259568 308898 259610 309134
rect 259846 308898 259888 309134
rect 259568 308866 259888 308898
rect 290288 309454 290608 309486
rect 290288 309218 290330 309454
rect 290566 309218 290608 309454
rect 290288 309134 290608 309218
rect 290288 308898 290330 309134
rect 290566 308898 290608 309134
rect 290288 308866 290608 308898
rect 321008 309454 321328 309486
rect 321008 309218 321050 309454
rect 321286 309218 321328 309454
rect 321008 309134 321328 309218
rect 321008 308898 321050 309134
rect 321286 308898 321328 309134
rect 321008 308866 321328 308898
rect 351728 309454 352048 309486
rect 351728 309218 351770 309454
rect 352006 309218 352048 309454
rect 351728 309134 352048 309218
rect 351728 308898 351770 309134
rect 352006 308898 352048 309134
rect 351728 308866 352048 308898
rect 382448 309454 382768 309486
rect 382448 309218 382490 309454
rect 382726 309218 382768 309454
rect 382448 309134 382768 309218
rect 382448 308898 382490 309134
rect 382726 308898 382768 309134
rect 382448 308866 382768 308898
rect 413168 309454 413488 309486
rect 413168 309218 413210 309454
rect 413446 309218 413488 309454
rect 413168 309134 413488 309218
rect 413168 308898 413210 309134
rect 413446 308898 413488 309134
rect 413168 308866 413488 308898
rect 443888 309454 444208 309486
rect 443888 309218 443930 309454
rect 444166 309218 444208 309454
rect 443888 309134 444208 309218
rect 443888 308898 443930 309134
rect 444166 308898 444208 309134
rect 443888 308866 444208 308898
rect 474608 309454 474928 309486
rect 474608 309218 474650 309454
rect 474886 309218 474928 309454
rect 474608 309134 474928 309218
rect 474608 308898 474650 309134
rect 474886 308898 474928 309134
rect 474608 308866 474928 308898
rect 505328 309454 505648 309486
rect 505328 309218 505370 309454
rect 505606 309218 505648 309454
rect 505328 309134 505648 309218
rect 505328 308898 505370 309134
rect 505606 308898 505648 309134
rect 505328 308866 505648 308898
rect 536048 309454 536368 309486
rect 536048 309218 536090 309454
rect 536326 309218 536368 309454
rect 536048 309134 536368 309218
rect 536048 308898 536090 309134
rect 536326 308898 536368 309134
rect 536048 308866 536368 308898
rect 244208 291454 244528 291486
rect 244208 291218 244250 291454
rect 244486 291218 244528 291454
rect 244208 291134 244528 291218
rect 244208 290898 244250 291134
rect 244486 290898 244528 291134
rect 244208 290866 244528 290898
rect 274928 291454 275248 291486
rect 274928 291218 274970 291454
rect 275206 291218 275248 291454
rect 274928 291134 275248 291218
rect 274928 290898 274970 291134
rect 275206 290898 275248 291134
rect 274928 290866 275248 290898
rect 305648 291454 305968 291486
rect 305648 291218 305690 291454
rect 305926 291218 305968 291454
rect 305648 291134 305968 291218
rect 305648 290898 305690 291134
rect 305926 290898 305968 291134
rect 305648 290866 305968 290898
rect 336368 291454 336688 291486
rect 336368 291218 336410 291454
rect 336646 291218 336688 291454
rect 336368 291134 336688 291218
rect 336368 290898 336410 291134
rect 336646 290898 336688 291134
rect 336368 290866 336688 290898
rect 367088 291454 367408 291486
rect 367088 291218 367130 291454
rect 367366 291218 367408 291454
rect 367088 291134 367408 291218
rect 367088 290898 367130 291134
rect 367366 290898 367408 291134
rect 367088 290866 367408 290898
rect 397808 291454 398128 291486
rect 397808 291218 397850 291454
rect 398086 291218 398128 291454
rect 397808 291134 398128 291218
rect 397808 290898 397850 291134
rect 398086 290898 398128 291134
rect 397808 290866 398128 290898
rect 428528 291454 428848 291486
rect 428528 291218 428570 291454
rect 428806 291218 428848 291454
rect 428528 291134 428848 291218
rect 428528 290898 428570 291134
rect 428806 290898 428848 291134
rect 428528 290866 428848 290898
rect 459248 291454 459568 291486
rect 459248 291218 459290 291454
rect 459526 291218 459568 291454
rect 459248 291134 459568 291218
rect 459248 290898 459290 291134
rect 459526 290898 459568 291134
rect 459248 290866 459568 290898
rect 489968 291454 490288 291486
rect 489968 291218 490010 291454
rect 490246 291218 490288 291454
rect 489968 291134 490288 291218
rect 489968 290898 490010 291134
rect 490246 290898 490288 291134
rect 489968 290866 490288 290898
rect 520688 291454 521008 291486
rect 520688 291218 520730 291454
rect 520966 291218 521008 291454
rect 520688 291134 521008 291218
rect 520688 290898 520730 291134
rect 520966 290898 521008 291134
rect 520688 290866 521008 290898
rect 259568 273454 259888 273486
rect 259568 273218 259610 273454
rect 259846 273218 259888 273454
rect 259568 273134 259888 273218
rect 259568 272898 259610 273134
rect 259846 272898 259888 273134
rect 259568 272866 259888 272898
rect 290288 273454 290608 273486
rect 290288 273218 290330 273454
rect 290566 273218 290608 273454
rect 290288 273134 290608 273218
rect 290288 272898 290330 273134
rect 290566 272898 290608 273134
rect 290288 272866 290608 272898
rect 321008 273454 321328 273486
rect 321008 273218 321050 273454
rect 321286 273218 321328 273454
rect 321008 273134 321328 273218
rect 321008 272898 321050 273134
rect 321286 272898 321328 273134
rect 321008 272866 321328 272898
rect 351728 273454 352048 273486
rect 351728 273218 351770 273454
rect 352006 273218 352048 273454
rect 351728 273134 352048 273218
rect 351728 272898 351770 273134
rect 352006 272898 352048 273134
rect 351728 272866 352048 272898
rect 382448 273454 382768 273486
rect 382448 273218 382490 273454
rect 382726 273218 382768 273454
rect 382448 273134 382768 273218
rect 382448 272898 382490 273134
rect 382726 272898 382768 273134
rect 382448 272866 382768 272898
rect 413168 273454 413488 273486
rect 413168 273218 413210 273454
rect 413446 273218 413488 273454
rect 413168 273134 413488 273218
rect 413168 272898 413210 273134
rect 413446 272898 413488 273134
rect 413168 272866 413488 272898
rect 443888 273454 444208 273486
rect 443888 273218 443930 273454
rect 444166 273218 444208 273454
rect 443888 273134 444208 273218
rect 443888 272898 443930 273134
rect 444166 272898 444208 273134
rect 443888 272866 444208 272898
rect 474608 273454 474928 273486
rect 474608 273218 474650 273454
rect 474886 273218 474928 273454
rect 474608 273134 474928 273218
rect 474608 272898 474650 273134
rect 474886 272898 474928 273134
rect 474608 272866 474928 272898
rect 505328 273454 505648 273486
rect 505328 273218 505370 273454
rect 505606 273218 505648 273454
rect 505328 273134 505648 273218
rect 505328 272898 505370 273134
rect 505606 272898 505648 273134
rect 505328 272866 505648 272898
rect 536048 273454 536368 273486
rect 536048 273218 536090 273454
rect 536326 273218 536368 273454
rect 536048 273134 536368 273218
rect 536048 272898 536090 273134
rect 536326 272898 536368 273134
rect 536048 272866 536368 272898
rect 244208 255454 244528 255486
rect 244208 255218 244250 255454
rect 244486 255218 244528 255454
rect 244208 255134 244528 255218
rect 244208 254898 244250 255134
rect 244486 254898 244528 255134
rect 244208 254866 244528 254898
rect 274928 255454 275248 255486
rect 274928 255218 274970 255454
rect 275206 255218 275248 255454
rect 274928 255134 275248 255218
rect 274928 254898 274970 255134
rect 275206 254898 275248 255134
rect 274928 254866 275248 254898
rect 305648 255454 305968 255486
rect 305648 255218 305690 255454
rect 305926 255218 305968 255454
rect 305648 255134 305968 255218
rect 305648 254898 305690 255134
rect 305926 254898 305968 255134
rect 305648 254866 305968 254898
rect 336368 255454 336688 255486
rect 336368 255218 336410 255454
rect 336646 255218 336688 255454
rect 336368 255134 336688 255218
rect 336368 254898 336410 255134
rect 336646 254898 336688 255134
rect 336368 254866 336688 254898
rect 367088 255454 367408 255486
rect 367088 255218 367130 255454
rect 367366 255218 367408 255454
rect 367088 255134 367408 255218
rect 367088 254898 367130 255134
rect 367366 254898 367408 255134
rect 367088 254866 367408 254898
rect 397808 255454 398128 255486
rect 397808 255218 397850 255454
rect 398086 255218 398128 255454
rect 397808 255134 398128 255218
rect 397808 254898 397850 255134
rect 398086 254898 398128 255134
rect 397808 254866 398128 254898
rect 428528 255454 428848 255486
rect 428528 255218 428570 255454
rect 428806 255218 428848 255454
rect 428528 255134 428848 255218
rect 428528 254898 428570 255134
rect 428806 254898 428848 255134
rect 428528 254866 428848 254898
rect 459248 255454 459568 255486
rect 459248 255218 459290 255454
rect 459526 255218 459568 255454
rect 459248 255134 459568 255218
rect 459248 254898 459290 255134
rect 459526 254898 459568 255134
rect 459248 254866 459568 254898
rect 489968 255454 490288 255486
rect 489968 255218 490010 255454
rect 490246 255218 490288 255454
rect 489968 255134 490288 255218
rect 489968 254898 490010 255134
rect 490246 254898 490288 255134
rect 489968 254866 490288 254898
rect 520688 255454 521008 255486
rect 520688 255218 520730 255454
rect 520966 255218 521008 255454
rect 520688 255134 521008 255218
rect 520688 254898 520730 255134
rect 520966 254898 521008 255134
rect 520688 254866 521008 254898
rect 259568 237454 259888 237486
rect 259568 237218 259610 237454
rect 259846 237218 259888 237454
rect 259568 237134 259888 237218
rect 259568 236898 259610 237134
rect 259846 236898 259888 237134
rect 259568 236866 259888 236898
rect 290288 237454 290608 237486
rect 290288 237218 290330 237454
rect 290566 237218 290608 237454
rect 290288 237134 290608 237218
rect 290288 236898 290330 237134
rect 290566 236898 290608 237134
rect 290288 236866 290608 236898
rect 321008 237454 321328 237486
rect 321008 237218 321050 237454
rect 321286 237218 321328 237454
rect 321008 237134 321328 237218
rect 321008 236898 321050 237134
rect 321286 236898 321328 237134
rect 321008 236866 321328 236898
rect 351728 237454 352048 237486
rect 351728 237218 351770 237454
rect 352006 237218 352048 237454
rect 351728 237134 352048 237218
rect 351728 236898 351770 237134
rect 352006 236898 352048 237134
rect 351728 236866 352048 236898
rect 382448 237454 382768 237486
rect 382448 237218 382490 237454
rect 382726 237218 382768 237454
rect 382448 237134 382768 237218
rect 382448 236898 382490 237134
rect 382726 236898 382768 237134
rect 382448 236866 382768 236898
rect 413168 237454 413488 237486
rect 413168 237218 413210 237454
rect 413446 237218 413488 237454
rect 413168 237134 413488 237218
rect 413168 236898 413210 237134
rect 413446 236898 413488 237134
rect 413168 236866 413488 236898
rect 443888 237454 444208 237486
rect 443888 237218 443930 237454
rect 444166 237218 444208 237454
rect 443888 237134 444208 237218
rect 443888 236898 443930 237134
rect 444166 236898 444208 237134
rect 443888 236866 444208 236898
rect 474608 237454 474928 237486
rect 474608 237218 474650 237454
rect 474886 237218 474928 237454
rect 474608 237134 474928 237218
rect 474608 236898 474650 237134
rect 474886 236898 474928 237134
rect 474608 236866 474928 236898
rect 505328 237454 505648 237486
rect 505328 237218 505370 237454
rect 505606 237218 505648 237454
rect 505328 237134 505648 237218
rect 505328 236898 505370 237134
rect 505606 236898 505648 237134
rect 505328 236866 505648 236898
rect 536048 237454 536368 237486
rect 536048 237218 536090 237454
rect 536326 237218 536368 237454
rect 536048 237134 536368 237218
rect 536048 236898 536090 237134
rect 536326 236898 536368 237134
rect 536048 236866 536368 236898
rect 244208 219454 244528 219486
rect 244208 219218 244250 219454
rect 244486 219218 244528 219454
rect 244208 219134 244528 219218
rect 244208 218898 244250 219134
rect 244486 218898 244528 219134
rect 244208 218866 244528 218898
rect 274928 219454 275248 219486
rect 274928 219218 274970 219454
rect 275206 219218 275248 219454
rect 274928 219134 275248 219218
rect 274928 218898 274970 219134
rect 275206 218898 275248 219134
rect 274928 218866 275248 218898
rect 305648 219454 305968 219486
rect 305648 219218 305690 219454
rect 305926 219218 305968 219454
rect 305648 219134 305968 219218
rect 305648 218898 305690 219134
rect 305926 218898 305968 219134
rect 305648 218866 305968 218898
rect 336368 219454 336688 219486
rect 336368 219218 336410 219454
rect 336646 219218 336688 219454
rect 336368 219134 336688 219218
rect 336368 218898 336410 219134
rect 336646 218898 336688 219134
rect 336368 218866 336688 218898
rect 367088 219454 367408 219486
rect 367088 219218 367130 219454
rect 367366 219218 367408 219454
rect 367088 219134 367408 219218
rect 367088 218898 367130 219134
rect 367366 218898 367408 219134
rect 367088 218866 367408 218898
rect 397808 219454 398128 219486
rect 397808 219218 397850 219454
rect 398086 219218 398128 219454
rect 397808 219134 398128 219218
rect 397808 218898 397850 219134
rect 398086 218898 398128 219134
rect 397808 218866 398128 218898
rect 428528 219454 428848 219486
rect 428528 219218 428570 219454
rect 428806 219218 428848 219454
rect 428528 219134 428848 219218
rect 428528 218898 428570 219134
rect 428806 218898 428848 219134
rect 428528 218866 428848 218898
rect 459248 219454 459568 219486
rect 459248 219218 459290 219454
rect 459526 219218 459568 219454
rect 459248 219134 459568 219218
rect 459248 218898 459290 219134
rect 459526 218898 459568 219134
rect 459248 218866 459568 218898
rect 489968 219454 490288 219486
rect 489968 219218 490010 219454
rect 490246 219218 490288 219454
rect 489968 219134 490288 219218
rect 489968 218898 490010 219134
rect 490246 218898 490288 219134
rect 489968 218866 490288 218898
rect 520688 219454 521008 219486
rect 520688 219218 520730 219454
rect 520966 219218 521008 219454
rect 520688 219134 521008 219218
rect 520688 218898 520730 219134
rect 520966 218898 521008 219134
rect 520688 218866 521008 218898
rect 259568 201454 259888 201486
rect 259568 201218 259610 201454
rect 259846 201218 259888 201454
rect 259568 201134 259888 201218
rect 259568 200898 259610 201134
rect 259846 200898 259888 201134
rect 259568 200866 259888 200898
rect 290288 201454 290608 201486
rect 290288 201218 290330 201454
rect 290566 201218 290608 201454
rect 290288 201134 290608 201218
rect 290288 200898 290330 201134
rect 290566 200898 290608 201134
rect 290288 200866 290608 200898
rect 321008 201454 321328 201486
rect 321008 201218 321050 201454
rect 321286 201218 321328 201454
rect 321008 201134 321328 201218
rect 321008 200898 321050 201134
rect 321286 200898 321328 201134
rect 321008 200866 321328 200898
rect 351728 201454 352048 201486
rect 351728 201218 351770 201454
rect 352006 201218 352048 201454
rect 351728 201134 352048 201218
rect 351728 200898 351770 201134
rect 352006 200898 352048 201134
rect 351728 200866 352048 200898
rect 382448 201454 382768 201486
rect 382448 201218 382490 201454
rect 382726 201218 382768 201454
rect 382448 201134 382768 201218
rect 382448 200898 382490 201134
rect 382726 200898 382768 201134
rect 382448 200866 382768 200898
rect 413168 201454 413488 201486
rect 413168 201218 413210 201454
rect 413446 201218 413488 201454
rect 413168 201134 413488 201218
rect 413168 200898 413210 201134
rect 413446 200898 413488 201134
rect 413168 200866 413488 200898
rect 443888 201454 444208 201486
rect 443888 201218 443930 201454
rect 444166 201218 444208 201454
rect 443888 201134 444208 201218
rect 443888 200898 443930 201134
rect 444166 200898 444208 201134
rect 443888 200866 444208 200898
rect 474608 201454 474928 201486
rect 474608 201218 474650 201454
rect 474886 201218 474928 201454
rect 474608 201134 474928 201218
rect 474608 200898 474650 201134
rect 474886 200898 474928 201134
rect 474608 200866 474928 200898
rect 505328 201454 505648 201486
rect 505328 201218 505370 201454
rect 505606 201218 505648 201454
rect 505328 201134 505648 201218
rect 505328 200898 505370 201134
rect 505606 200898 505648 201134
rect 505328 200866 505648 200898
rect 536048 201454 536368 201486
rect 536048 201218 536090 201454
rect 536326 201218 536368 201454
rect 536048 201134 536368 201218
rect 536048 200898 536090 201134
rect 536326 200898 536368 201134
rect 536048 200866 536368 200898
rect 244208 183454 244528 183486
rect 244208 183218 244250 183454
rect 244486 183218 244528 183454
rect 244208 183134 244528 183218
rect 244208 182898 244250 183134
rect 244486 182898 244528 183134
rect 244208 182866 244528 182898
rect 274928 183454 275248 183486
rect 274928 183218 274970 183454
rect 275206 183218 275248 183454
rect 274928 183134 275248 183218
rect 274928 182898 274970 183134
rect 275206 182898 275248 183134
rect 274928 182866 275248 182898
rect 305648 183454 305968 183486
rect 305648 183218 305690 183454
rect 305926 183218 305968 183454
rect 305648 183134 305968 183218
rect 305648 182898 305690 183134
rect 305926 182898 305968 183134
rect 305648 182866 305968 182898
rect 336368 183454 336688 183486
rect 336368 183218 336410 183454
rect 336646 183218 336688 183454
rect 336368 183134 336688 183218
rect 336368 182898 336410 183134
rect 336646 182898 336688 183134
rect 336368 182866 336688 182898
rect 367088 183454 367408 183486
rect 367088 183218 367130 183454
rect 367366 183218 367408 183454
rect 367088 183134 367408 183218
rect 367088 182898 367130 183134
rect 367366 182898 367408 183134
rect 367088 182866 367408 182898
rect 397808 183454 398128 183486
rect 397808 183218 397850 183454
rect 398086 183218 398128 183454
rect 397808 183134 398128 183218
rect 397808 182898 397850 183134
rect 398086 182898 398128 183134
rect 397808 182866 398128 182898
rect 428528 183454 428848 183486
rect 428528 183218 428570 183454
rect 428806 183218 428848 183454
rect 428528 183134 428848 183218
rect 428528 182898 428570 183134
rect 428806 182898 428848 183134
rect 428528 182866 428848 182898
rect 459248 183454 459568 183486
rect 459248 183218 459290 183454
rect 459526 183218 459568 183454
rect 459248 183134 459568 183218
rect 459248 182898 459290 183134
rect 459526 182898 459568 183134
rect 459248 182866 459568 182898
rect 489968 183454 490288 183486
rect 489968 183218 490010 183454
rect 490246 183218 490288 183454
rect 489968 183134 490288 183218
rect 489968 182898 490010 183134
rect 490246 182898 490288 183134
rect 489968 182866 490288 182898
rect 520688 183454 521008 183486
rect 520688 183218 520730 183454
rect 520966 183218 521008 183454
rect 520688 183134 521008 183218
rect 520688 182898 520730 183134
rect 520966 182898 521008 183134
rect 520688 182866 521008 182898
rect 536790 179757 536850 596803
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 482000 542414 506898
rect 545514 691174 546134 706202
rect 545514 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 546134 691174
rect 545514 690854 546134 690938
rect 545514 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 546134 690854
rect 545514 655174 546134 690618
rect 545514 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 546134 655174
rect 545514 654854 546134 654938
rect 545514 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 546134 654854
rect 545514 619174 546134 654618
rect 545514 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 546134 619174
rect 545514 618854 546134 618938
rect 545514 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 546134 618854
rect 545514 583174 546134 618618
rect 545514 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 546134 583174
rect 545514 582854 546134 582938
rect 545514 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 546134 582854
rect 545514 547174 546134 582618
rect 545514 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 546134 547174
rect 545514 546854 546134 546938
rect 545514 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 546134 546854
rect 545514 511174 546134 546618
rect 545514 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 546134 511174
rect 545514 510854 546134 510938
rect 545514 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 546134 510854
rect 545514 475174 546134 510618
rect 545514 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 546134 475174
rect 545514 474854 546134 474938
rect 545514 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 546134 474854
rect 545514 439174 546134 474618
rect 545514 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 546134 439174
rect 545514 438854 546134 438938
rect 545514 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 546134 438854
rect 545514 403174 546134 438618
rect 545514 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 546134 403174
rect 545514 402854 546134 402938
rect 545514 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 546134 402854
rect 545514 367174 546134 402618
rect 545514 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 546134 367174
rect 545514 366854 546134 366938
rect 545514 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 546134 366854
rect 545514 331174 546134 366618
rect 545514 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 546134 331174
rect 545514 330854 546134 330938
rect 545514 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 546134 330854
rect 545514 295174 546134 330618
rect 545514 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 546134 295174
rect 545514 294854 546134 294938
rect 545514 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 546134 294854
rect 545514 259174 546134 294618
rect 545514 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 546134 259174
rect 545514 258854 546134 258938
rect 545514 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 546134 258854
rect 545514 223174 546134 258618
rect 545514 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 546134 223174
rect 545514 222854 546134 222938
rect 545514 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 546134 222854
rect 545514 187174 546134 222618
rect 545514 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 546134 187174
rect 545514 186854 546134 186938
rect 545514 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 546134 186854
rect 536787 179756 536853 179757
rect 536787 179692 536788 179756
rect 536852 179692 536853 179756
rect 536787 179691 536853 179692
rect 239259 178940 239325 178941
rect 239259 178876 239260 178940
rect 239324 178876 239325 178940
rect 239259 178875 239325 178876
rect 235794 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 236414 165454
rect 235794 165134 236414 165218
rect 235794 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 236414 165134
rect 235794 129454 236414 164898
rect 235794 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 236414 129454
rect 235794 129134 236414 129218
rect 235794 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 236414 129134
rect 235794 93454 236414 128898
rect 235794 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 236414 93454
rect 235794 93134 236414 93218
rect 235794 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 236414 93134
rect 235794 57454 236414 92898
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -1306 236414 20898
rect 235794 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 236414 -1306
rect 235794 -1626 236414 -1542
rect 235794 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 236414 -1626
rect 235794 -1894 236414 -1862
rect 239514 169174 240134 178000
rect 239514 168938 239546 169174
rect 239782 168938 239866 169174
rect 240102 168938 240134 169174
rect 239514 168854 240134 168938
rect 239514 168618 239546 168854
rect 239782 168618 239866 168854
rect 240102 168618 240134 168854
rect 239514 133174 240134 168618
rect 239514 132938 239546 133174
rect 239782 132938 239866 133174
rect 240102 132938 240134 133174
rect 239514 132854 240134 132938
rect 239514 132618 239546 132854
rect 239782 132618 239866 132854
rect 240102 132618 240134 132854
rect 239514 97174 240134 132618
rect 239514 96938 239546 97174
rect 239782 96938 239866 97174
rect 240102 96938 240134 97174
rect 239514 96854 240134 96938
rect 239514 96618 239546 96854
rect 239782 96618 239866 96854
rect 240102 96618 240134 96854
rect 239514 61174 240134 96618
rect 239514 60938 239546 61174
rect 239782 60938 239866 61174
rect 240102 60938 240134 61174
rect 239514 60854 240134 60938
rect 239514 60618 239546 60854
rect 239782 60618 239866 60854
rect 240102 60618 240134 60854
rect 239514 25174 240134 60618
rect 239514 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 240134 25174
rect 239514 24854 240134 24938
rect 239514 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 240134 24854
rect 239514 -3226 240134 24618
rect 239514 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 240134 -3226
rect 239514 -3546 240134 -3462
rect 239514 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 240134 -3546
rect 239514 -3814 240134 -3782
rect 243234 172894 243854 178000
rect 243234 172658 243266 172894
rect 243502 172658 243586 172894
rect 243822 172658 243854 172894
rect 243234 172574 243854 172658
rect 243234 172338 243266 172574
rect 243502 172338 243586 172574
rect 243822 172338 243854 172574
rect 243234 136894 243854 172338
rect 243234 136658 243266 136894
rect 243502 136658 243586 136894
rect 243822 136658 243854 136894
rect 243234 136574 243854 136658
rect 243234 136338 243266 136574
rect 243502 136338 243586 136574
rect 243822 136338 243854 136574
rect 243234 100894 243854 136338
rect 243234 100658 243266 100894
rect 243502 100658 243586 100894
rect 243822 100658 243854 100894
rect 243234 100574 243854 100658
rect 243234 100338 243266 100574
rect 243502 100338 243586 100574
rect 243822 100338 243854 100574
rect 243234 64894 243854 100338
rect 243234 64658 243266 64894
rect 243502 64658 243586 64894
rect 243822 64658 243854 64894
rect 243234 64574 243854 64658
rect 243234 64338 243266 64574
rect 243502 64338 243586 64574
rect 243822 64338 243854 64574
rect 243234 28894 243854 64338
rect 243234 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 243854 28894
rect 243234 28574 243854 28658
rect 243234 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 243854 28574
rect 243234 -5146 243854 28338
rect 243234 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 243854 -5146
rect 243234 -5466 243854 -5382
rect 243234 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 243854 -5466
rect 243234 -5734 243854 -5702
rect 246954 176614 247574 178000
rect 246954 176378 246986 176614
rect 247222 176378 247306 176614
rect 247542 176378 247574 176614
rect 246954 176294 247574 176378
rect 246954 176058 246986 176294
rect 247222 176058 247306 176294
rect 247542 176058 247574 176294
rect 246954 140614 247574 176058
rect 246954 140378 246986 140614
rect 247222 140378 247306 140614
rect 247542 140378 247574 140614
rect 246954 140294 247574 140378
rect 246954 140058 246986 140294
rect 247222 140058 247306 140294
rect 247542 140058 247574 140294
rect 246954 104614 247574 140058
rect 246954 104378 246986 104614
rect 247222 104378 247306 104614
rect 247542 104378 247574 104614
rect 246954 104294 247574 104378
rect 246954 104058 246986 104294
rect 247222 104058 247306 104294
rect 247542 104058 247574 104294
rect 246954 68614 247574 104058
rect 246954 68378 246986 68614
rect 247222 68378 247306 68614
rect 247542 68378 247574 68614
rect 246954 68294 247574 68378
rect 246954 68058 246986 68294
rect 247222 68058 247306 68294
rect 247542 68058 247574 68294
rect 246954 32614 247574 68058
rect 246954 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 247574 32614
rect 246954 32294 247574 32378
rect 246954 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 247574 32294
rect 228954 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 229574 -6106
rect 228954 -6426 229574 -6342
rect 228954 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 229574 -6426
rect 228954 -7654 229574 -6662
rect 246954 -7066 247574 32058
rect 253794 147454 254414 178000
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 253794 111454 254414 146898
rect 253794 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 254414 111454
rect 253794 111134 254414 111218
rect 253794 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 254414 111134
rect 253794 75454 254414 110898
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -1894 254414 -902
rect 257514 151174 258134 178000
rect 257514 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 258134 151174
rect 257514 150854 258134 150938
rect 257514 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 258134 150854
rect 257514 115174 258134 150618
rect 257514 114938 257546 115174
rect 257782 114938 257866 115174
rect 258102 114938 258134 115174
rect 257514 114854 258134 114938
rect 257514 114618 257546 114854
rect 257782 114618 257866 114854
rect 258102 114618 258134 114854
rect 257514 79174 258134 114618
rect 257514 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 258134 79174
rect 257514 78854 258134 78938
rect 257514 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 258134 78854
rect 257514 43174 258134 78618
rect 257514 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 258134 43174
rect 257514 42854 258134 42938
rect 257514 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 258134 42854
rect 257514 7174 258134 42618
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 257514 -2266 258134 6618
rect 257514 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 258134 -2266
rect 257514 -2586 258134 -2502
rect 257514 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 258134 -2586
rect 257514 -3814 258134 -2822
rect 261234 154894 261854 178000
rect 261234 154658 261266 154894
rect 261502 154658 261586 154894
rect 261822 154658 261854 154894
rect 261234 154574 261854 154658
rect 261234 154338 261266 154574
rect 261502 154338 261586 154574
rect 261822 154338 261854 154574
rect 261234 118894 261854 154338
rect 261234 118658 261266 118894
rect 261502 118658 261586 118894
rect 261822 118658 261854 118894
rect 261234 118574 261854 118658
rect 261234 118338 261266 118574
rect 261502 118338 261586 118574
rect 261822 118338 261854 118574
rect 261234 82894 261854 118338
rect 261234 82658 261266 82894
rect 261502 82658 261586 82894
rect 261822 82658 261854 82894
rect 261234 82574 261854 82658
rect 261234 82338 261266 82574
rect 261502 82338 261586 82574
rect 261822 82338 261854 82574
rect 261234 46894 261854 82338
rect 261234 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 261854 46894
rect 261234 46574 261854 46658
rect 261234 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 261854 46574
rect 261234 10894 261854 46338
rect 261234 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 261854 10894
rect 261234 10574 261854 10658
rect 261234 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 261854 10574
rect 261234 -4186 261854 10338
rect 261234 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 261854 -4186
rect 261234 -4506 261854 -4422
rect 261234 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 261854 -4506
rect 261234 -5734 261854 -4742
rect 264954 158614 265574 178000
rect 264954 158378 264986 158614
rect 265222 158378 265306 158614
rect 265542 158378 265574 158614
rect 264954 158294 265574 158378
rect 264954 158058 264986 158294
rect 265222 158058 265306 158294
rect 265542 158058 265574 158294
rect 264954 122614 265574 158058
rect 264954 122378 264986 122614
rect 265222 122378 265306 122614
rect 265542 122378 265574 122614
rect 264954 122294 265574 122378
rect 264954 122058 264986 122294
rect 265222 122058 265306 122294
rect 265542 122058 265574 122294
rect 264954 86614 265574 122058
rect 264954 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 265574 86614
rect 264954 86294 265574 86378
rect 264954 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 265574 86294
rect 264954 50614 265574 86058
rect 264954 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 265574 50614
rect 264954 50294 265574 50378
rect 264954 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 265574 50294
rect 264954 14614 265574 50058
rect 264954 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 265574 14614
rect 264954 14294 265574 14378
rect 264954 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 265574 14294
rect 246954 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 247574 -7066
rect 246954 -7386 247574 -7302
rect 246954 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 247574 -7386
rect 246954 -7654 247574 -7622
rect 264954 -6106 265574 14058
rect 271794 165454 272414 178000
rect 271794 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 272414 165454
rect 271794 165134 272414 165218
rect 271794 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 272414 165134
rect 271794 129454 272414 164898
rect 271794 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 272414 129454
rect 271794 129134 272414 129218
rect 271794 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 272414 129134
rect 271794 93454 272414 128898
rect 271794 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 272414 93454
rect 271794 93134 272414 93218
rect 271794 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 272414 93134
rect 271794 57454 272414 92898
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -1306 272414 20898
rect 271794 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 272414 -1306
rect 271794 -1626 272414 -1542
rect 271794 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 272414 -1626
rect 271794 -1894 272414 -1862
rect 275514 169174 276134 178000
rect 275514 168938 275546 169174
rect 275782 168938 275866 169174
rect 276102 168938 276134 169174
rect 275514 168854 276134 168938
rect 275514 168618 275546 168854
rect 275782 168618 275866 168854
rect 276102 168618 276134 168854
rect 275514 133174 276134 168618
rect 275514 132938 275546 133174
rect 275782 132938 275866 133174
rect 276102 132938 276134 133174
rect 275514 132854 276134 132938
rect 275514 132618 275546 132854
rect 275782 132618 275866 132854
rect 276102 132618 276134 132854
rect 275514 97174 276134 132618
rect 275514 96938 275546 97174
rect 275782 96938 275866 97174
rect 276102 96938 276134 97174
rect 275514 96854 276134 96938
rect 275514 96618 275546 96854
rect 275782 96618 275866 96854
rect 276102 96618 276134 96854
rect 275514 61174 276134 96618
rect 275514 60938 275546 61174
rect 275782 60938 275866 61174
rect 276102 60938 276134 61174
rect 275514 60854 276134 60938
rect 275514 60618 275546 60854
rect 275782 60618 275866 60854
rect 276102 60618 276134 60854
rect 275514 25174 276134 60618
rect 275514 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 276134 25174
rect 275514 24854 276134 24938
rect 275514 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 276134 24854
rect 275514 -3226 276134 24618
rect 275514 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 276134 -3226
rect 275514 -3546 276134 -3462
rect 275514 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 276134 -3546
rect 275514 -3814 276134 -3782
rect 279234 172894 279854 178000
rect 279234 172658 279266 172894
rect 279502 172658 279586 172894
rect 279822 172658 279854 172894
rect 279234 172574 279854 172658
rect 279234 172338 279266 172574
rect 279502 172338 279586 172574
rect 279822 172338 279854 172574
rect 279234 136894 279854 172338
rect 279234 136658 279266 136894
rect 279502 136658 279586 136894
rect 279822 136658 279854 136894
rect 279234 136574 279854 136658
rect 279234 136338 279266 136574
rect 279502 136338 279586 136574
rect 279822 136338 279854 136574
rect 279234 100894 279854 136338
rect 279234 100658 279266 100894
rect 279502 100658 279586 100894
rect 279822 100658 279854 100894
rect 279234 100574 279854 100658
rect 279234 100338 279266 100574
rect 279502 100338 279586 100574
rect 279822 100338 279854 100574
rect 279234 64894 279854 100338
rect 279234 64658 279266 64894
rect 279502 64658 279586 64894
rect 279822 64658 279854 64894
rect 279234 64574 279854 64658
rect 279234 64338 279266 64574
rect 279502 64338 279586 64574
rect 279822 64338 279854 64574
rect 279234 28894 279854 64338
rect 279234 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 279854 28894
rect 279234 28574 279854 28658
rect 279234 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 279854 28574
rect 279234 -5146 279854 28338
rect 279234 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 279854 -5146
rect 279234 -5466 279854 -5382
rect 279234 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 279854 -5466
rect 279234 -5734 279854 -5702
rect 282954 176614 283574 178000
rect 282954 176378 282986 176614
rect 283222 176378 283306 176614
rect 283542 176378 283574 176614
rect 282954 176294 283574 176378
rect 282954 176058 282986 176294
rect 283222 176058 283306 176294
rect 283542 176058 283574 176294
rect 282954 140614 283574 176058
rect 282954 140378 282986 140614
rect 283222 140378 283306 140614
rect 283542 140378 283574 140614
rect 282954 140294 283574 140378
rect 282954 140058 282986 140294
rect 283222 140058 283306 140294
rect 283542 140058 283574 140294
rect 282954 104614 283574 140058
rect 282954 104378 282986 104614
rect 283222 104378 283306 104614
rect 283542 104378 283574 104614
rect 282954 104294 283574 104378
rect 282954 104058 282986 104294
rect 283222 104058 283306 104294
rect 283542 104058 283574 104294
rect 282954 68614 283574 104058
rect 282954 68378 282986 68614
rect 283222 68378 283306 68614
rect 283542 68378 283574 68614
rect 282954 68294 283574 68378
rect 282954 68058 282986 68294
rect 283222 68058 283306 68294
rect 283542 68058 283574 68294
rect 282954 32614 283574 68058
rect 282954 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 283574 32614
rect 282954 32294 283574 32378
rect 282954 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 283574 32294
rect 264954 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 265574 -6106
rect 264954 -6426 265574 -6342
rect 264954 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 265574 -6426
rect 264954 -7654 265574 -6662
rect 282954 -7066 283574 32058
rect 289794 147454 290414 178000
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 289794 111454 290414 146898
rect 289794 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 290414 111454
rect 289794 111134 290414 111218
rect 289794 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 290414 111134
rect 289794 75454 290414 110898
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -1894 290414 -902
rect 293514 151174 294134 178000
rect 293514 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 294134 151174
rect 293514 150854 294134 150938
rect 293514 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 294134 150854
rect 293514 115174 294134 150618
rect 293514 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 294134 115174
rect 293514 114854 294134 114938
rect 293514 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 294134 114854
rect 293514 79174 294134 114618
rect 293514 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 294134 79174
rect 293514 78854 294134 78938
rect 293514 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 294134 78854
rect 293514 43174 294134 78618
rect 293514 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 294134 43174
rect 293514 42854 294134 42938
rect 293514 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 294134 42854
rect 293514 7174 294134 42618
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 293514 -2266 294134 6618
rect 293514 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 294134 -2266
rect 293514 -2586 294134 -2502
rect 293514 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 294134 -2586
rect 293514 -3814 294134 -2822
rect 297234 154894 297854 178000
rect 297234 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 297854 154894
rect 297234 154574 297854 154658
rect 297234 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 297854 154574
rect 297234 118894 297854 154338
rect 297234 118658 297266 118894
rect 297502 118658 297586 118894
rect 297822 118658 297854 118894
rect 297234 118574 297854 118658
rect 297234 118338 297266 118574
rect 297502 118338 297586 118574
rect 297822 118338 297854 118574
rect 297234 82894 297854 118338
rect 297234 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 297854 82894
rect 297234 82574 297854 82658
rect 297234 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 297854 82574
rect 297234 46894 297854 82338
rect 297234 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 297854 46894
rect 297234 46574 297854 46658
rect 297234 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 297854 46574
rect 297234 10894 297854 46338
rect 297234 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 297854 10894
rect 297234 10574 297854 10658
rect 297234 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 297854 10574
rect 297234 -4186 297854 10338
rect 297234 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 297854 -4186
rect 297234 -4506 297854 -4422
rect 297234 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 297854 -4506
rect 297234 -5734 297854 -4742
rect 300954 158614 301574 178000
rect 300954 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 301574 158614
rect 300954 158294 301574 158378
rect 300954 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 301574 158294
rect 300954 122614 301574 158058
rect 300954 122378 300986 122614
rect 301222 122378 301306 122614
rect 301542 122378 301574 122614
rect 300954 122294 301574 122378
rect 300954 122058 300986 122294
rect 301222 122058 301306 122294
rect 301542 122058 301574 122294
rect 300954 86614 301574 122058
rect 300954 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 301574 86614
rect 300954 86294 301574 86378
rect 300954 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 301574 86294
rect 300954 50614 301574 86058
rect 300954 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 301574 50614
rect 300954 50294 301574 50378
rect 300954 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 301574 50294
rect 300954 14614 301574 50058
rect 300954 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 301574 14614
rect 300954 14294 301574 14378
rect 300954 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 301574 14294
rect 282954 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 283574 -7066
rect 282954 -7386 283574 -7302
rect 282954 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 283574 -7386
rect 282954 -7654 283574 -7622
rect 300954 -6106 301574 14058
rect 307794 165454 308414 178000
rect 307794 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 308414 165454
rect 307794 165134 308414 165218
rect 307794 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 308414 165134
rect 307794 129454 308414 164898
rect 307794 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 308414 129454
rect 307794 129134 308414 129218
rect 307794 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 308414 129134
rect 307794 93454 308414 128898
rect 307794 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 308414 93454
rect 307794 93134 308414 93218
rect 307794 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 308414 93134
rect 307794 57454 308414 92898
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -1306 308414 20898
rect 307794 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 308414 -1306
rect 307794 -1626 308414 -1542
rect 307794 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 308414 -1626
rect 307794 -1894 308414 -1862
rect 311514 169174 312134 178000
rect 311514 168938 311546 169174
rect 311782 168938 311866 169174
rect 312102 168938 312134 169174
rect 311514 168854 312134 168938
rect 311514 168618 311546 168854
rect 311782 168618 311866 168854
rect 312102 168618 312134 168854
rect 311514 133174 312134 168618
rect 311514 132938 311546 133174
rect 311782 132938 311866 133174
rect 312102 132938 312134 133174
rect 311514 132854 312134 132938
rect 311514 132618 311546 132854
rect 311782 132618 311866 132854
rect 312102 132618 312134 132854
rect 311514 97174 312134 132618
rect 311514 96938 311546 97174
rect 311782 96938 311866 97174
rect 312102 96938 312134 97174
rect 311514 96854 312134 96938
rect 311514 96618 311546 96854
rect 311782 96618 311866 96854
rect 312102 96618 312134 96854
rect 311514 61174 312134 96618
rect 311514 60938 311546 61174
rect 311782 60938 311866 61174
rect 312102 60938 312134 61174
rect 311514 60854 312134 60938
rect 311514 60618 311546 60854
rect 311782 60618 311866 60854
rect 312102 60618 312134 60854
rect 311514 25174 312134 60618
rect 311514 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 312134 25174
rect 311514 24854 312134 24938
rect 311514 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 312134 24854
rect 311514 -3226 312134 24618
rect 311514 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 312134 -3226
rect 311514 -3546 312134 -3462
rect 311514 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 312134 -3546
rect 311514 -3814 312134 -3782
rect 315234 172894 315854 178000
rect 315234 172658 315266 172894
rect 315502 172658 315586 172894
rect 315822 172658 315854 172894
rect 315234 172574 315854 172658
rect 315234 172338 315266 172574
rect 315502 172338 315586 172574
rect 315822 172338 315854 172574
rect 315234 136894 315854 172338
rect 315234 136658 315266 136894
rect 315502 136658 315586 136894
rect 315822 136658 315854 136894
rect 315234 136574 315854 136658
rect 315234 136338 315266 136574
rect 315502 136338 315586 136574
rect 315822 136338 315854 136574
rect 315234 100894 315854 136338
rect 315234 100658 315266 100894
rect 315502 100658 315586 100894
rect 315822 100658 315854 100894
rect 315234 100574 315854 100658
rect 315234 100338 315266 100574
rect 315502 100338 315586 100574
rect 315822 100338 315854 100574
rect 315234 64894 315854 100338
rect 315234 64658 315266 64894
rect 315502 64658 315586 64894
rect 315822 64658 315854 64894
rect 315234 64574 315854 64658
rect 315234 64338 315266 64574
rect 315502 64338 315586 64574
rect 315822 64338 315854 64574
rect 315234 28894 315854 64338
rect 315234 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 315854 28894
rect 315234 28574 315854 28658
rect 315234 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 315854 28574
rect 315234 -5146 315854 28338
rect 315234 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 315854 -5146
rect 315234 -5466 315854 -5382
rect 315234 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 315854 -5466
rect 315234 -5734 315854 -5702
rect 318954 176614 319574 178000
rect 318954 176378 318986 176614
rect 319222 176378 319306 176614
rect 319542 176378 319574 176614
rect 318954 176294 319574 176378
rect 318954 176058 318986 176294
rect 319222 176058 319306 176294
rect 319542 176058 319574 176294
rect 318954 140614 319574 176058
rect 318954 140378 318986 140614
rect 319222 140378 319306 140614
rect 319542 140378 319574 140614
rect 318954 140294 319574 140378
rect 318954 140058 318986 140294
rect 319222 140058 319306 140294
rect 319542 140058 319574 140294
rect 318954 104614 319574 140058
rect 318954 104378 318986 104614
rect 319222 104378 319306 104614
rect 319542 104378 319574 104614
rect 318954 104294 319574 104378
rect 318954 104058 318986 104294
rect 319222 104058 319306 104294
rect 319542 104058 319574 104294
rect 318954 68614 319574 104058
rect 318954 68378 318986 68614
rect 319222 68378 319306 68614
rect 319542 68378 319574 68614
rect 318954 68294 319574 68378
rect 318954 68058 318986 68294
rect 319222 68058 319306 68294
rect 319542 68058 319574 68294
rect 318954 32614 319574 68058
rect 318954 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 319574 32614
rect 318954 32294 319574 32378
rect 318954 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 319574 32294
rect 300954 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 301574 -6106
rect 300954 -6426 301574 -6342
rect 300954 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 301574 -6426
rect 300954 -7654 301574 -6662
rect 318954 -7066 319574 32058
rect 325794 147454 326414 178000
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 325794 111454 326414 146898
rect 325794 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 326414 111454
rect 325794 111134 326414 111218
rect 325794 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 326414 111134
rect 325794 75454 326414 110898
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -1894 326414 -902
rect 329514 151174 330134 178000
rect 329514 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 330134 151174
rect 329514 150854 330134 150938
rect 329514 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 330134 150854
rect 329514 115174 330134 150618
rect 329514 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 330134 115174
rect 329514 114854 330134 114938
rect 329514 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 330134 114854
rect 329514 79174 330134 114618
rect 329514 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 330134 79174
rect 329514 78854 330134 78938
rect 329514 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 330134 78854
rect 329514 43174 330134 78618
rect 329514 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 330134 43174
rect 329514 42854 330134 42938
rect 329514 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 330134 42854
rect 329514 7174 330134 42618
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -2266 330134 6618
rect 329514 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 330134 -2266
rect 329514 -2586 330134 -2502
rect 329514 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 330134 -2586
rect 329514 -3814 330134 -2822
rect 333234 154894 333854 178000
rect 333234 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 333854 154894
rect 333234 154574 333854 154658
rect 333234 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 333854 154574
rect 333234 118894 333854 154338
rect 333234 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 333854 118894
rect 333234 118574 333854 118658
rect 333234 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 333854 118574
rect 333234 82894 333854 118338
rect 333234 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 333854 82894
rect 333234 82574 333854 82658
rect 333234 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 333854 82574
rect 333234 46894 333854 82338
rect 333234 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 333854 46894
rect 333234 46574 333854 46658
rect 333234 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 333854 46574
rect 333234 10894 333854 46338
rect 333234 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 333854 10894
rect 333234 10574 333854 10658
rect 333234 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 333854 10574
rect 333234 -4186 333854 10338
rect 333234 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 333854 -4186
rect 333234 -4506 333854 -4422
rect 333234 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 333854 -4506
rect 333234 -5734 333854 -4742
rect 336954 158614 337574 178000
rect 336954 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 337574 158614
rect 336954 158294 337574 158378
rect 336954 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 337574 158294
rect 336954 122614 337574 158058
rect 336954 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 337574 122614
rect 336954 122294 337574 122378
rect 336954 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 337574 122294
rect 336954 86614 337574 122058
rect 336954 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 337574 86614
rect 336954 86294 337574 86378
rect 336954 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 337574 86294
rect 336954 50614 337574 86058
rect 336954 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 337574 50614
rect 336954 50294 337574 50378
rect 336954 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 337574 50294
rect 336954 14614 337574 50058
rect 336954 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 337574 14614
rect 336954 14294 337574 14378
rect 336954 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 337574 14294
rect 318954 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 319574 -7066
rect 318954 -7386 319574 -7302
rect 318954 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 319574 -7386
rect 318954 -7654 319574 -7622
rect 336954 -6106 337574 14058
rect 343794 165454 344414 178000
rect 343794 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 344414 165454
rect 343794 165134 344414 165218
rect 343794 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 344414 165134
rect 343794 129454 344414 164898
rect 343794 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 344414 129454
rect 343794 129134 344414 129218
rect 343794 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 344414 129134
rect 343794 93454 344414 128898
rect 343794 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 344414 93454
rect 343794 93134 344414 93218
rect 343794 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 344414 93134
rect 343794 57454 344414 92898
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -1306 344414 20898
rect 343794 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 344414 -1306
rect 343794 -1626 344414 -1542
rect 343794 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 344414 -1626
rect 343794 -1894 344414 -1862
rect 347514 169174 348134 178000
rect 347514 168938 347546 169174
rect 347782 168938 347866 169174
rect 348102 168938 348134 169174
rect 347514 168854 348134 168938
rect 347514 168618 347546 168854
rect 347782 168618 347866 168854
rect 348102 168618 348134 168854
rect 347514 133174 348134 168618
rect 347514 132938 347546 133174
rect 347782 132938 347866 133174
rect 348102 132938 348134 133174
rect 347514 132854 348134 132938
rect 347514 132618 347546 132854
rect 347782 132618 347866 132854
rect 348102 132618 348134 132854
rect 347514 97174 348134 132618
rect 347514 96938 347546 97174
rect 347782 96938 347866 97174
rect 348102 96938 348134 97174
rect 347514 96854 348134 96938
rect 347514 96618 347546 96854
rect 347782 96618 347866 96854
rect 348102 96618 348134 96854
rect 347514 61174 348134 96618
rect 347514 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 348134 61174
rect 347514 60854 348134 60938
rect 347514 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 348134 60854
rect 347514 25174 348134 60618
rect 347514 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 348134 25174
rect 347514 24854 348134 24938
rect 347514 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 348134 24854
rect 347514 -3226 348134 24618
rect 347514 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 348134 -3226
rect 347514 -3546 348134 -3462
rect 347514 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 348134 -3546
rect 347514 -3814 348134 -3782
rect 351234 172894 351854 178000
rect 351234 172658 351266 172894
rect 351502 172658 351586 172894
rect 351822 172658 351854 172894
rect 351234 172574 351854 172658
rect 351234 172338 351266 172574
rect 351502 172338 351586 172574
rect 351822 172338 351854 172574
rect 351234 136894 351854 172338
rect 351234 136658 351266 136894
rect 351502 136658 351586 136894
rect 351822 136658 351854 136894
rect 351234 136574 351854 136658
rect 351234 136338 351266 136574
rect 351502 136338 351586 136574
rect 351822 136338 351854 136574
rect 351234 100894 351854 136338
rect 351234 100658 351266 100894
rect 351502 100658 351586 100894
rect 351822 100658 351854 100894
rect 351234 100574 351854 100658
rect 351234 100338 351266 100574
rect 351502 100338 351586 100574
rect 351822 100338 351854 100574
rect 351234 64894 351854 100338
rect 351234 64658 351266 64894
rect 351502 64658 351586 64894
rect 351822 64658 351854 64894
rect 351234 64574 351854 64658
rect 351234 64338 351266 64574
rect 351502 64338 351586 64574
rect 351822 64338 351854 64574
rect 351234 28894 351854 64338
rect 351234 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 351854 28894
rect 351234 28574 351854 28658
rect 351234 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 351854 28574
rect 351234 -5146 351854 28338
rect 351234 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 351854 -5146
rect 351234 -5466 351854 -5382
rect 351234 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 351854 -5466
rect 351234 -5734 351854 -5702
rect 354954 176614 355574 178000
rect 354954 176378 354986 176614
rect 355222 176378 355306 176614
rect 355542 176378 355574 176614
rect 354954 176294 355574 176378
rect 354954 176058 354986 176294
rect 355222 176058 355306 176294
rect 355542 176058 355574 176294
rect 354954 140614 355574 176058
rect 354954 140378 354986 140614
rect 355222 140378 355306 140614
rect 355542 140378 355574 140614
rect 354954 140294 355574 140378
rect 354954 140058 354986 140294
rect 355222 140058 355306 140294
rect 355542 140058 355574 140294
rect 354954 104614 355574 140058
rect 354954 104378 354986 104614
rect 355222 104378 355306 104614
rect 355542 104378 355574 104614
rect 354954 104294 355574 104378
rect 354954 104058 354986 104294
rect 355222 104058 355306 104294
rect 355542 104058 355574 104294
rect 354954 68614 355574 104058
rect 354954 68378 354986 68614
rect 355222 68378 355306 68614
rect 355542 68378 355574 68614
rect 354954 68294 355574 68378
rect 354954 68058 354986 68294
rect 355222 68058 355306 68294
rect 355542 68058 355574 68294
rect 354954 32614 355574 68058
rect 354954 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 355574 32614
rect 354954 32294 355574 32378
rect 354954 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 355574 32294
rect 336954 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 337574 -6106
rect 336954 -6426 337574 -6342
rect 336954 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 337574 -6426
rect 336954 -7654 337574 -6662
rect 354954 -7066 355574 32058
rect 361794 147454 362414 178000
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -1894 362414 -902
rect 365514 151174 366134 178000
rect 365514 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 366134 151174
rect 365514 150854 366134 150938
rect 365514 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 366134 150854
rect 365514 115174 366134 150618
rect 365514 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 366134 115174
rect 365514 114854 366134 114938
rect 365514 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 366134 114854
rect 365514 79174 366134 114618
rect 365514 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 366134 79174
rect 365514 78854 366134 78938
rect 365514 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 366134 78854
rect 365514 43174 366134 78618
rect 365514 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 366134 43174
rect 365514 42854 366134 42938
rect 365514 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 366134 42854
rect 365514 7174 366134 42618
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 365514 -2266 366134 6618
rect 365514 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 366134 -2266
rect 365514 -2586 366134 -2502
rect 365514 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 366134 -2586
rect 365514 -3814 366134 -2822
rect 369234 154894 369854 178000
rect 369234 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 369854 154894
rect 369234 154574 369854 154658
rect 369234 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 369854 154574
rect 369234 118894 369854 154338
rect 369234 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 369854 118894
rect 369234 118574 369854 118658
rect 369234 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 369854 118574
rect 369234 82894 369854 118338
rect 369234 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 369854 82894
rect 369234 82574 369854 82658
rect 369234 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 369854 82574
rect 369234 46894 369854 82338
rect 369234 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 369854 46894
rect 369234 46574 369854 46658
rect 369234 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 369854 46574
rect 369234 10894 369854 46338
rect 369234 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 369854 10894
rect 369234 10574 369854 10658
rect 369234 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 369854 10574
rect 369234 -4186 369854 10338
rect 369234 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 369854 -4186
rect 369234 -4506 369854 -4422
rect 369234 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 369854 -4506
rect 369234 -5734 369854 -4742
rect 372954 158614 373574 178000
rect 372954 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 373574 158614
rect 372954 158294 373574 158378
rect 372954 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 373574 158294
rect 372954 122614 373574 158058
rect 372954 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 373574 122614
rect 372954 122294 373574 122378
rect 372954 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 373574 122294
rect 372954 86614 373574 122058
rect 372954 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 373574 86614
rect 372954 86294 373574 86378
rect 372954 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 373574 86294
rect 372954 50614 373574 86058
rect 372954 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 373574 50614
rect 372954 50294 373574 50378
rect 372954 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 373574 50294
rect 372954 14614 373574 50058
rect 372954 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 373574 14614
rect 372954 14294 373574 14378
rect 372954 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 373574 14294
rect 354954 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 355574 -7066
rect 354954 -7386 355574 -7302
rect 354954 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 355574 -7386
rect 354954 -7654 355574 -7622
rect 372954 -6106 373574 14058
rect 379794 165454 380414 178000
rect 379794 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 380414 165454
rect 379794 165134 380414 165218
rect 379794 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 380414 165134
rect 379794 129454 380414 164898
rect 379794 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 380414 129454
rect 379794 129134 380414 129218
rect 379794 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 380414 129134
rect 379794 93454 380414 128898
rect 379794 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 380414 93454
rect 379794 93134 380414 93218
rect 379794 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 380414 93134
rect 379794 57454 380414 92898
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -1306 380414 20898
rect 379794 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 380414 -1306
rect 379794 -1626 380414 -1542
rect 379794 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 380414 -1626
rect 379794 -1894 380414 -1862
rect 383514 169174 384134 178000
rect 383514 168938 383546 169174
rect 383782 168938 383866 169174
rect 384102 168938 384134 169174
rect 383514 168854 384134 168938
rect 383514 168618 383546 168854
rect 383782 168618 383866 168854
rect 384102 168618 384134 168854
rect 383514 133174 384134 168618
rect 383514 132938 383546 133174
rect 383782 132938 383866 133174
rect 384102 132938 384134 133174
rect 383514 132854 384134 132938
rect 383514 132618 383546 132854
rect 383782 132618 383866 132854
rect 384102 132618 384134 132854
rect 383514 97174 384134 132618
rect 383514 96938 383546 97174
rect 383782 96938 383866 97174
rect 384102 96938 384134 97174
rect 383514 96854 384134 96938
rect 383514 96618 383546 96854
rect 383782 96618 383866 96854
rect 384102 96618 384134 96854
rect 383514 61174 384134 96618
rect 383514 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 384134 61174
rect 383514 60854 384134 60938
rect 383514 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 384134 60854
rect 383514 25174 384134 60618
rect 383514 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 384134 25174
rect 383514 24854 384134 24938
rect 383514 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 384134 24854
rect 383514 -3226 384134 24618
rect 383514 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 384134 -3226
rect 383514 -3546 384134 -3462
rect 383514 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 384134 -3546
rect 383514 -3814 384134 -3782
rect 387234 172894 387854 178000
rect 387234 172658 387266 172894
rect 387502 172658 387586 172894
rect 387822 172658 387854 172894
rect 387234 172574 387854 172658
rect 387234 172338 387266 172574
rect 387502 172338 387586 172574
rect 387822 172338 387854 172574
rect 387234 136894 387854 172338
rect 387234 136658 387266 136894
rect 387502 136658 387586 136894
rect 387822 136658 387854 136894
rect 387234 136574 387854 136658
rect 387234 136338 387266 136574
rect 387502 136338 387586 136574
rect 387822 136338 387854 136574
rect 387234 100894 387854 136338
rect 387234 100658 387266 100894
rect 387502 100658 387586 100894
rect 387822 100658 387854 100894
rect 387234 100574 387854 100658
rect 387234 100338 387266 100574
rect 387502 100338 387586 100574
rect 387822 100338 387854 100574
rect 387234 64894 387854 100338
rect 387234 64658 387266 64894
rect 387502 64658 387586 64894
rect 387822 64658 387854 64894
rect 387234 64574 387854 64658
rect 387234 64338 387266 64574
rect 387502 64338 387586 64574
rect 387822 64338 387854 64574
rect 387234 28894 387854 64338
rect 387234 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 387854 28894
rect 387234 28574 387854 28658
rect 387234 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 387854 28574
rect 387234 -5146 387854 28338
rect 387234 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 387854 -5146
rect 387234 -5466 387854 -5382
rect 387234 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 387854 -5466
rect 387234 -5734 387854 -5702
rect 390954 176614 391574 178000
rect 390954 176378 390986 176614
rect 391222 176378 391306 176614
rect 391542 176378 391574 176614
rect 390954 176294 391574 176378
rect 390954 176058 390986 176294
rect 391222 176058 391306 176294
rect 391542 176058 391574 176294
rect 390954 140614 391574 176058
rect 390954 140378 390986 140614
rect 391222 140378 391306 140614
rect 391542 140378 391574 140614
rect 390954 140294 391574 140378
rect 390954 140058 390986 140294
rect 391222 140058 391306 140294
rect 391542 140058 391574 140294
rect 390954 104614 391574 140058
rect 390954 104378 390986 104614
rect 391222 104378 391306 104614
rect 391542 104378 391574 104614
rect 390954 104294 391574 104378
rect 390954 104058 390986 104294
rect 391222 104058 391306 104294
rect 391542 104058 391574 104294
rect 390954 68614 391574 104058
rect 390954 68378 390986 68614
rect 391222 68378 391306 68614
rect 391542 68378 391574 68614
rect 390954 68294 391574 68378
rect 390954 68058 390986 68294
rect 391222 68058 391306 68294
rect 391542 68058 391574 68294
rect 390954 32614 391574 68058
rect 390954 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 391574 32614
rect 390954 32294 391574 32378
rect 390954 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 391574 32294
rect 372954 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 373574 -6106
rect 372954 -6426 373574 -6342
rect 372954 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 373574 -6426
rect 372954 -7654 373574 -6662
rect 390954 -7066 391574 32058
rect 397794 147454 398414 178000
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -1894 398414 -902
rect 401514 151174 402134 178000
rect 401514 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 402134 151174
rect 401514 150854 402134 150938
rect 401514 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 402134 150854
rect 401514 115174 402134 150618
rect 401514 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 402134 115174
rect 401514 114854 402134 114938
rect 401514 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 402134 114854
rect 401514 79174 402134 114618
rect 401514 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 402134 79174
rect 401514 78854 402134 78938
rect 401514 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 402134 78854
rect 401514 43174 402134 78618
rect 401514 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 402134 43174
rect 401514 42854 402134 42938
rect 401514 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 402134 42854
rect 401514 7174 402134 42618
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -2266 402134 6618
rect 401514 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 402134 -2266
rect 401514 -2586 402134 -2502
rect 401514 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 402134 -2586
rect 401514 -3814 402134 -2822
rect 405234 154894 405854 178000
rect 405234 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 405854 154894
rect 405234 154574 405854 154658
rect 405234 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 405854 154574
rect 405234 118894 405854 154338
rect 405234 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 405854 118894
rect 405234 118574 405854 118658
rect 405234 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 405854 118574
rect 405234 82894 405854 118338
rect 405234 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 405854 82894
rect 405234 82574 405854 82658
rect 405234 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 405854 82574
rect 405234 46894 405854 82338
rect 405234 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 405854 46894
rect 405234 46574 405854 46658
rect 405234 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 405854 46574
rect 405234 10894 405854 46338
rect 405234 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 405854 10894
rect 405234 10574 405854 10658
rect 405234 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 405854 10574
rect 405234 -4186 405854 10338
rect 405234 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 405854 -4186
rect 405234 -4506 405854 -4422
rect 405234 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 405854 -4506
rect 405234 -5734 405854 -4742
rect 408954 158614 409574 178000
rect 408954 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 409574 158614
rect 408954 158294 409574 158378
rect 408954 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 409574 158294
rect 408954 122614 409574 158058
rect 408954 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 409574 122614
rect 408954 122294 409574 122378
rect 408954 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 409574 122294
rect 408954 86614 409574 122058
rect 408954 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 409574 86614
rect 408954 86294 409574 86378
rect 408954 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 409574 86294
rect 408954 50614 409574 86058
rect 408954 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 409574 50614
rect 408954 50294 409574 50378
rect 408954 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 409574 50294
rect 408954 14614 409574 50058
rect 408954 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 409574 14614
rect 408954 14294 409574 14378
rect 408954 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 409574 14294
rect 390954 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 391574 -7066
rect 390954 -7386 391574 -7302
rect 390954 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 391574 -7386
rect 390954 -7654 391574 -7622
rect 408954 -6106 409574 14058
rect 415794 165454 416414 178000
rect 415794 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 416414 165454
rect 415794 165134 416414 165218
rect 415794 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 416414 165134
rect 415794 129454 416414 164898
rect 415794 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 416414 129454
rect 415794 129134 416414 129218
rect 415794 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 416414 129134
rect 415794 93454 416414 128898
rect 415794 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 416414 93454
rect 415794 93134 416414 93218
rect 415794 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 416414 93134
rect 415794 57454 416414 92898
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -1306 416414 20898
rect 415794 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 416414 -1306
rect 415794 -1626 416414 -1542
rect 415794 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 416414 -1626
rect 415794 -1894 416414 -1862
rect 419514 169174 420134 178000
rect 419514 168938 419546 169174
rect 419782 168938 419866 169174
rect 420102 168938 420134 169174
rect 419514 168854 420134 168938
rect 419514 168618 419546 168854
rect 419782 168618 419866 168854
rect 420102 168618 420134 168854
rect 419514 133174 420134 168618
rect 419514 132938 419546 133174
rect 419782 132938 419866 133174
rect 420102 132938 420134 133174
rect 419514 132854 420134 132938
rect 419514 132618 419546 132854
rect 419782 132618 419866 132854
rect 420102 132618 420134 132854
rect 419514 97174 420134 132618
rect 419514 96938 419546 97174
rect 419782 96938 419866 97174
rect 420102 96938 420134 97174
rect 419514 96854 420134 96938
rect 419514 96618 419546 96854
rect 419782 96618 419866 96854
rect 420102 96618 420134 96854
rect 419514 61174 420134 96618
rect 419514 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 420134 61174
rect 419514 60854 420134 60938
rect 419514 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 420134 60854
rect 419514 25174 420134 60618
rect 419514 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 420134 25174
rect 419514 24854 420134 24938
rect 419514 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 420134 24854
rect 419514 -3226 420134 24618
rect 419514 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 420134 -3226
rect 419514 -3546 420134 -3462
rect 419514 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 420134 -3546
rect 419514 -3814 420134 -3782
rect 423234 172894 423854 178000
rect 423234 172658 423266 172894
rect 423502 172658 423586 172894
rect 423822 172658 423854 172894
rect 423234 172574 423854 172658
rect 423234 172338 423266 172574
rect 423502 172338 423586 172574
rect 423822 172338 423854 172574
rect 423234 136894 423854 172338
rect 423234 136658 423266 136894
rect 423502 136658 423586 136894
rect 423822 136658 423854 136894
rect 423234 136574 423854 136658
rect 423234 136338 423266 136574
rect 423502 136338 423586 136574
rect 423822 136338 423854 136574
rect 423234 100894 423854 136338
rect 423234 100658 423266 100894
rect 423502 100658 423586 100894
rect 423822 100658 423854 100894
rect 423234 100574 423854 100658
rect 423234 100338 423266 100574
rect 423502 100338 423586 100574
rect 423822 100338 423854 100574
rect 423234 64894 423854 100338
rect 423234 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 423854 64894
rect 423234 64574 423854 64658
rect 423234 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 423854 64574
rect 423234 28894 423854 64338
rect 423234 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 423854 28894
rect 423234 28574 423854 28658
rect 423234 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 423854 28574
rect 423234 -5146 423854 28338
rect 423234 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 423854 -5146
rect 423234 -5466 423854 -5382
rect 423234 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 423854 -5466
rect 423234 -5734 423854 -5702
rect 426954 176614 427574 178000
rect 426954 176378 426986 176614
rect 427222 176378 427306 176614
rect 427542 176378 427574 176614
rect 426954 176294 427574 176378
rect 426954 176058 426986 176294
rect 427222 176058 427306 176294
rect 427542 176058 427574 176294
rect 426954 140614 427574 176058
rect 426954 140378 426986 140614
rect 427222 140378 427306 140614
rect 427542 140378 427574 140614
rect 426954 140294 427574 140378
rect 426954 140058 426986 140294
rect 427222 140058 427306 140294
rect 427542 140058 427574 140294
rect 426954 104614 427574 140058
rect 426954 104378 426986 104614
rect 427222 104378 427306 104614
rect 427542 104378 427574 104614
rect 426954 104294 427574 104378
rect 426954 104058 426986 104294
rect 427222 104058 427306 104294
rect 427542 104058 427574 104294
rect 426954 68614 427574 104058
rect 426954 68378 426986 68614
rect 427222 68378 427306 68614
rect 427542 68378 427574 68614
rect 426954 68294 427574 68378
rect 426954 68058 426986 68294
rect 427222 68058 427306 68294
rect 427542 68058 427574 68294
rect 426954 32614 427574 68058
rect 426954 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 427574 32614
rect 426954 32294 427574 32378
rect 426954 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 427574 32294
rect 408954 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 409574 -6106
rect 408954 -6426 409574 -6342
rect 408954 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 409574 -6426
rect 408954 -7654 409574 -6662
rect 426954 -7066 427574 32058
rect 433794 147454 434414 178000
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 111454 434414 146898
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -1894 434414 -902
rect 437514 151174 438134 178000
rect 437514 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 438134 151174
rect 437514 150854 438134 150938
rect 437514 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 438134 150854
rect 437514 115174 438134 150618
rect 437514 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 438134 115174
rect 437514 114854 438134 114938
rect 437514 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 438134 114854
rect 437514 79174 438134 114618
rect 437514 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 438134 79174
rect 437514 78854 438134 78938
rect 437514 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 438134 78854
rect 437514 43174 438134 78618
rect 437514 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 438134 43174
rect 437514 42854 438134 42938
rect 437514 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 438134 42854
rect 437514 7174 438134 42618
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -2266 438134 6618
rect 437514 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 438134 -2266
rect 437514 -2586 438134 -2502
rect 437514 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 438134 -2586
rect 437514 -3814 438134 -2822
rect 441234 154894 441854 178000
rect 441234 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 441854 154894
rect 441234 154574 441854 154658
rect 441234 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 441854 154574
rect 441234 118894 441854 154338
rect 441234 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 441854 118894
rect 441234 118574 441854 118658
rect 441234 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 441854 118574
rect 441234 82894 441854 118338
rect 441234 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 441854 82894
rect 441234 82574 441854 82658
rect 441234 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 441854 82574
rect 441234 46894 441854 82338
rect 441234 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 441854 46894
rect 441234 46574 441854 46658
rect 441234 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 441854 46574
rect 441234 10894 441854 46338
rect 441234 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 441854 10894
rect 441234 10574 441854 10658
rect 441234 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 441854 10574
rect 441234 -4186 441854 10338
rect 441234 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 441854 -4186
rect 441234 -4506 441854 -4422
rect 441234 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 441854 -4506
rect 441234 -5734 441854 -4742
rect 444954 158614 445574 178000
rect 444954 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 445574 158614
rect 444954 158294 445574 158378
rect 444954 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 445574 158294
rect 444954 122614 445574 158058
rect 444954 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 445574 122614
rect 444954 122294 445574 122378
rect 444954 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 445574 122294
rect 444954 86614 445574 122058
rect 444954 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 445574 86614
rect 444954 86294 445574 86378
rect 444954 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 445574 86294
rect 444954 50614 445574 86058
rect 444954 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 445574 50614
rect 444954 50294 445574 50378
rect 444954 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 445574 50294
rect 444954 14614 445574 50058
rect 444954 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 445574 14614
rect 444954 14294 445574 14378
rect 444954 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 445574 14294
rect 426954 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 427574 -7066
rect 426954 -7386 427574 -7302
rect 426954 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 427574 -7386
rect 426954 -7654 427574 -7622
rect 444954 -6106 445574 14058
rect 451794 165454 452414 178000
rect 451794 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 452414 165454
rect 451794 165134 452414 165218
rect 451794 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 452414 165134
rect 451794 129454 452414 164898
rect 451794 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 452414 129454
rect 451794 129134 452414 129218
rect 451794 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 452414 129134
rect 451794 93454 452414 128898
rect 451794 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 452414 93454
rect 451794 93134 452414 93218
rect 451794 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 452414 93134
rect 451794 57454 452414 92898
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -1306 452414 20898
rect 451794 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 452414 -1306
rect 451794 -1626 452414 -1542
rect 451794 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 452414 -1626
rect 451794 -1894 452414 -1862
rect 455514 169174 456134 178000
rect 455514 168938 455546 169174
rect 455782 168938 455866 169174
rect 456102 168938 456134 169174
rect 455514 168854 456134 168938
rect 455514 168618 455546 168854
rect 455782 168618 455866 168854
rect 456102 168618 456134 168854
rect 455514 133174 456134 168618
rect 455514 132938 455546 133174
rect 455782 132938 455866 133174
rect 456102 132938 456134 133174
rect 455514 132854 456134 132938
rect 455514 132618 455546 132854
rect 455782 132618 455866 132854
rect 456102 132618 456134 132854
rect 455514 97174 456134 132618
rect 455514 96938 455546 97174
rect 455782 96938 455866 97174
rect 456102 96938 456134 97174
rect 455514 96854 456134 96938
rect 455514 96618 455546 96854
rect 455782 96618 455866 96854
rect 456102 96618 456134 96854
rect 455514 61174 456134 96618
rect 455514 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 456134 61174
rect 455514 60854 456134 60938
rect 455514 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 456134 60854
rect 455514 25174 456134 60618
rect 455514 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 456134 25174
rect 455514 24854 456134 24938
rect 455514 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 456134 24854
rect 455514 -3226 456134 24618
rect 455514 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 456134 -3226
rect 455514 -3546 456134 -3462
rect 455514 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 456134 -3546
rect 455514 -3814 456134 -3782
rect 459234 172894 459854 178000
rect 459234 172658 459266 172894
rect 459502 172658 459586 172894
rect 459822 172658 459854 172894
rect 459234 172574 459854 172658
rect 459234 172338 459266 172574
rect 459502 172338 459586 172574
rect 459822 172338 459854 172574
rect 459234 136894 459854 172338
rect 459234 136658 459266 136894
rect 459502 136658 459586 136894
rect 459822 136658 459854 136894
rect 459234 136574 459854 136658
rect 459234 136338 459266 136574
rect 459502 136338 459586 136574
rect 459822 136338 459854 136574
rect 459234 100894 459854 136338
rect 459234 100658 459266 100894
rect 459502 100658 459586 100894
rect 459822 100658 459854 100894
rect 459234 100574 459854 100658
rect 459234 100338 459266 100574
rect 459502 100338 459586 100574
rect 459822 100338 459854 100574
rect 459234 64894 459854 100338
rect 459234 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 459854 64894
rect 459234 64574 459854 64658
rect 459234 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 459854 64574
rect 459234 28894 459854 64338
rect 459234 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 459854 28894
rect 459234 28574 459854 28658
rect 459234 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 459854 28574
rect 459234 -5146 459854 28338
rect 459234 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 459854 -5146
rect 459234 -5466 459854 -5382
rect 459234 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 459854 -5466
rect 459234 -5734 459854 -5702
rect 462954 176614 463574 178000
rect 462954 176378 462986 176614
rect 463222 176378 463306 176614
rect 463542 176378 463574 176614
rect 462954 176294 463574 176378
rect 462954 176058 462986 176294
rect 463222 176058 463306 176294
rect 463542 176058 463574 176294
rect 462954 140614 463574 176058
rect 462954 140378 462986 140614
rect 463222 140378 463306 140614
rect 463542 140378 463574 140614
rect 462954 140294 463574 140378
rect 462954 140058 462986 140294
rect 463222 140058 463306 140294
rect 463542 140058 463574 140294
rect 462954 104614 463574 140058
rect 462954 104378 462986 104614
rect 463222 104378 463306 104614
rect 463542 104378 463574 104614
rect 462954 104294 463574 104378
rect 462954 104058 462986 104294
rect 463222 104058 463306 104294
rect 463542 104058 463574 104294
rect 462954 68614 463574 104058
rect 462954 68378 462986 68614
rect 463222 68378 463306 68614
rect 463542 68378 463574 68614
rect 462954 68294 463574 68378
rect 462954 68058 462986 68294
rect 463222 68058 463306 68294
rect 463542 68058 463574 68294
rect 462954 32614 463574 68058
rect 462954 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 463574 32614
rect 462954 32294 463574 32378
rect 462954 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 463574 32294
rect 444954 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 445574 -6106
rect 444954 -6426 445574 -6342
rect 444954 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 445574 -6426
rect 444954 -7654 445574 -6662
rect 462954 -7066 463574 32058
rect 469794 147454 470414 178000
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -1894 470414 -902
rect 473514 151174 474134 178000
rect 473514 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 474134 151174
rect 473514 150854 474134 150938
rect 473514 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 474134 150854
rect 473514 115174 474134 150618
rect 473514 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 474134 115174
rect 473514 114854 474134 114938
rect 473514 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 474134 114854
rect 473514 79174 474134 114618
rect 473514 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 474134 79174
rect 473514 78854 474134 78938
rect 473514 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 474134 78854
rect 473514 43174 474134 78618
rect 473514 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 474134 43174
rect 473514 42854 474134 42938
rect 473514 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 474134 42854
rect 473514 7174 474134 42618
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -2266 474134 6618
rect 473514 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 474134 -2266
rect 473514 -2586 474134 -2502
rect 473514 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 474134 -2586
rect 473514 -3814 474134 -2822
rect 477234 154894 477854 178000
rect 477234 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 477854 154894
rect 477234 154574 477854 154658
rect 477234 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 477854 154574
rect 477234 118894 477854 154338
rect 477234 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 477854 118894
rect 477234 118574 477854 118658
rect 477234 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 477854 118574
rect 477234 82894 477854 118338
rect 477234 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 477854 82894
rect 477234 82574 477854 82658
rect 477234 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 477854 82574
rect 477234 46894 477854 82338
rect 477234 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 477854 46894
rect 477234 46574 477854 46658
rect 477234 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 477854 46574
rect 477234 10894 477854 46338
rect 477234 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 477854 10894
rect 477234 10574 477854 10658
rect 477234 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 477854 10574
rect 477234 -4186 477854 10338
rect 477234 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 477854 -4186
rect 477234 -4506 477854 -4422
rect 477234 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 477854 -4506
rect 477234 -5734 477854 -4742
rect 480954 158614 481574 178000
rect 480954 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 481574 158614
rect 480954 158294 481574 158378
rect 480954 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 481574 158294
rect 480954 122614 481574 158058
rect 480954 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 481574 122614
rect 480954 122294 481574 122378
rect 480954 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 481574 122294
rect 480954 86614 481574 122058
rect 480954 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 481574 86614
rect 480954 86294 481574 86378
rect 480954 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 481574 86294
rect 480954 50614 481574 86058
rect 480954 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 481574 50614
rect 480954 50294 481574 50378
rect 480954 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 481574 50294
rect 480954 14614 481574 50058
rect 480954 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 481574 14614
rect 480954 14294 481574 14378
rect 480954 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 481574 14294
rect 462954 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 463574 -7066
rect 462954 -7386 463574 -7302
rect 462954 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 463574 -7386
rect 462954 -7654 463574 -7622
rect 480954 -6106 481574 14058
rect 487794 165454 488414 178000
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 129454 488414 164898
rect 487794 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 488414 129454
rect 487794 129134 488414 129218
rect 487794 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 488414 129134
rect 487794 93454 488414 128898
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -1306 488414 20898
rect 487794 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 488414 -1306
rect 487794 -1626 488414 -1542
rect 487794 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 488414 -1626
rect 487794 -1894 488414 -1862
rect 491514 169174 492134 178000
rect 491514 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 492134 169174
rect 491514 168854 492134 168938
rect 491514 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 492134 168854
rect 491514 133174 492134 168618
rect 491514 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 492134 133174
rect 491514 132854 492134 132938
rect 491514 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 492134 132854
rect 491514 97174 492134 132618
rect 491514 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 492134 97174
rect 491514 96854 492134 96938
rect 491514 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 492134 96854
rect 491514 61174 492134 96618
rect 491514 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 492134 61174
rect 491514 60854 492134 60938
rect 491514 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 492134 60854
rect 491514 25174 492134 60618
rect 491514 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 492134 25174
rect 491514 24854 492134 24938
rect 491514 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 492134 24854
rect 491514 -3226 492134 24618
rect 491514 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 492134 -3226
rect 491514 -3546 492134 -3462
rect 491514 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 492134 -3546
rect 491514 -3814 492134 -3782
rect 495234 172894 495854 178000
rect 495234 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 495854 172894
rect 495234 172574 495854 172658
rect 495234 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 495854 172574
rect 495234 136894 495854 172338
rect 495234 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 495854 136894
rect 495234 136574 495854 136658
rect 495234 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 495854 136574
rect 495234 100894 495854 136338
rect 495234 100658 495266 100894
rect 495502 100658 495586 100894
rect 495822 100658 495854 100894
rect 495234 100574 495854 100658
rect 495234 100338 495266 100574
rect 495502 100338 495586 100574
rect 495822 100338 495854 100574
rect 495234 64894 495854 100338
rect 495234 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 495854 64894
rect 495234 64574 495854 64658
rect 495234 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 495854 64574
rect 495234 28894 495854 64338
rect 495234 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 495854 28894
rect 495234 28574 495854 28658
rect 495234 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 495854 28574
rect 495234 -5146 495854 28338
rect 495234 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 495854 -5146
rect 495234 -5466 495854 -5382
rect 495234 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 495854 -5466
rect 495234 -5734 495854 -5702
rect 498954 176614 499574 178000
rect 498954 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 499574 176614
rect 498954 176294 499574 176378
rect 498954 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 499574 176294
rect 498954 140614 499574 176058
rect 498954 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 499574 140614
rect 498954 140294 499574 140378
rect 498954 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 499574 140294
rect 498954 104614 499574 140058
rect 498954 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 499574 104614
rect 498954 104294 499574 104378
rect 498954 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 499574 104294
rect 498954 68614 499574 104058
rect 498954 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 499574 68614
rect 498954 68294 499574 68378
rect 498954 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 499574 68294
rect 498954 32614 499574 68058
rect 498954 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 499574 32614
rect 498954 32294 499574 32378
rect 498954 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 499574 32294
rect 480954 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 481574 -6106
rect 480954 -6426 481574 -6342
rect 480954 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 481574 -6426
rect 480954 -7654 481574 -6662
rect 498954 -7066 499574 32058
rect 505794 147454 506414 178000
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -1894 506414 -902
rect 509514 151174 510134 178000
rect 509514 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 510134 151174
rect 509514 150854 510134 150938
rect 509514 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 510134 150854
rect 509514 115174 510134 150618
rect 509514 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 510134 115174
rect 509514 114854 510134 114938
rect 509514 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 510134 114854
rect 509514 79174 510134 114618
rect 509514 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 510134 79174
rect 509514 78854 510134 78938
rect 509514 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 510134 78854
rect 509514 43174 510134 78618
rect 509514 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 510134 43174
rect 509514 42854 510134 42938
rect 509514 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 510134 42854
rect 509514 7174 510134 42618
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -2266 510134 6618
rect 509514 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 510134 -2266
rect 509514 -2586 510134 -2502
rect 509514 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 510134 -2586
rect 509514 -3814 510134 -2822
rect 513234 154894 513854 178000
rect 513234 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 513854 154894
rect 513234 154574 513854 154658
rect 513234 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 513854 154574
rect 513234 118894 513854 154338
rect 513234 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 513854 118894
rect 513234 118574 513854 118658
rect 513234 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 513854 118574
rect 513234 82894 513854 118338
rect 513234 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 513854 82894
rect 513234 82574 513854 82658
rect 513234 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 513854 82574
rect 513234 46894 513854 82338
rect 513234 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 513854 46894
rect 513234 46574 513854 46658
rect 513234 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 513854 46574
rect 513234 10894 513854 46338
rect 513234 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 513854 10894
rect 513234 10574 513854 10658
rect 513234 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 513854 10574
rect 513234 -4186 513854 10338
rect 513234 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 513854 -4186
rect 513234 -4506 513854 -4422
rect 513234 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 513854 -4506
rect 513234 -5734 513854 -4742
rect 516954 158614 517574 178000
rect 516954 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 517574 158614
rect 516954 158294 517574 158378
rect 516954 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 517574 158294
rect 516954 122614 517574 158058
rect 516954 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 517574 122614
rect 516954 122294 517574 122378
rect 516954 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 517574 122294
rect 516954 86614 517574 122058
rect 516954 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 517574 86614
rect 516954 86294 517574 86378
rect 516954 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 517574 86294
rect 516954 50614 517574 86058
rect 516954 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 517574 50614
rect 516954 50294 517574 50378
rect 516954 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 517574 50294
rect 516954 14614 517574 50058
rect 516954 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 517574 14614
rect 516954 14294 517574 14378
rect 516954 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 517574 14294
rect 498954 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 499574 -7066
rect 498954 -7386 499574 -7302
rect 498954 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 499574 -7386
rect 498954 -7654 499574 -7622
rect 516954 -6106 517574 14058
rect 523794 165454 524414 178000
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -1306 524414 20898
rect 523794 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 524414 -1306
rect 523794 -1626 524414 -1542
rect 523794 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 524414 -1626
rect 523794 -1894 524414 -1862
rect 527514 169174 528134 178000
rect 527514 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 528134 169174
rect 527514 168854 528134 168938
rect 527514 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 528134 168854
rect 527514 133174 528134 168618
rect 527514 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 528134 133174
rect 527514 132854 528134 132938
rect 527514 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 528134 132854
rect 527514 97174 528134 132618
rect 527514 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 528134 97174
rect 527514 96854 528134 96938
rect 527514 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 528134 96854
rect 527514 61174 528134 96618
rect 527514 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 528134 61174
rect 527514 60854 528134 60938
rect 527514 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 528134 60854
rect 527514 25174 528134 60618
rect 527514 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 528134 25174
rect 527514 24854 528134 24938
rect 527514 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 528134 24854
rect 527514 -3226 528134 24618
rect 527514 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 528134 -3226
rect 527514 -3546 528134 -3462
rect 527514 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 528134 -3546
rect 527514 -3814 528134 -3782
rect 531234 172894 531854 178000
rect 531234 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 531854 172894
rect 531234 172574 531854 172658
rect 531234 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 531854 172574
rect 531234 136894 531854 172338
rect 531234 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 531854 136894
rect 531234 136574 531854 136658
rect 531234 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 531854 136574
rect 531234 100894 531854 136338
rect 531234 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 531854 100894
rect 531234 100574 531854 100658
rect 531234 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 531854 100574
rect 531234 64894 531854 100338
rect 531234 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 531854 64894
rect 531234 64574 531854 64658
rect 531234 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 531854 64574
rect 531234 28894 531854 64338
rect 531234 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 531854 28894
rect 531234 28574 531854 28658
rect 531234 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 531854 28574
rect 531234 -5146 531854 28338
rect 531234 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 531854 -5146
rect 531234 -5466 531854 -5382
rect 531234 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 531854 -5466
rect 531234 -5734 531854 -5702
rect 534954 176614 535574 178000
rect 534954 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 535574 176614
rect 534954 176294 535574 176378
rect 534954 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 535574 176294
rect 534954 140614 535574 176058
rect 534954 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 535574 140614
rect 534954 140294 535574 140378
rect 534954 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 535574 140294
rect 534954 104614 535574 140058
rect 534954 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 535574 104614
rect 534954 104294 535574 104378
rect 534954 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 535574 104294
rect 534954 68614 535574 104058
rect 534954 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 535574 68614
rect 534954 68294 535574 68378
rect 534954 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 535574 68294
rect 534954 32614 535574 68058
rect 534954 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 535574 32614
rect 534954 32294 535574 32378
rect 534954 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 535574 32294
rect 516954 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 517574 -6106
rect 516954 -6426 517574 -6342
rect 516954 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 517574 -6426
rect 516954 -7654 517574 -6662
rect 534954 -7066 535574 32058
rect 541794 147454 542414 178000
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -1894 542414 -902
rect 545514 151174 546134 186618
rect 545514 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 546134 151174
rect 545514 150854 546134 150938
rect 545514 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 546134 150854
rect 545514 115174 546134 150618
rect 545514 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 546134 115174
rect 545514 114854 546134 114938
rect 545514 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 546134 114854
rect 545514 79174 546134 114618
rect 545514 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 546134 79174
rect 545514 78854 546134 78938
rect 545514 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 546134 78854
rect 545514 43174 546134 78618
rect 545514 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 546134 43174
rect 545514 42854 546134 42938
rect 545514 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 546134 42854
rect 545514 7174 546134 42618
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -2266 546134 6618
rect 545514 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 546134 -2266
rect 545514 -2586 546134 -2502
rect 545514 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 546134 -2586
rect 545514 -3814 546134 -2822
rect 549234 694894 549854 708122
rect 549234 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 549854 694894
rect 549234 694574 549854 694658
rect 549234 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 549854 694574
rect 549234 658894 549854 694338
rect 549234 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 549854 658894
rect 549234 658574 549854 658658
rect 549234 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 549854 658574
rect 549234 622894 549854 658338
rect 549234 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 549854 622894
rect 549234 622574 549854 622658
rect 549234 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 549854 622574
rect 549234 586894 549854 622338
rect 549234 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 549854 586894
rect 549234 586574 549854 586658
rect 549234 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 549854 586574
rect 549234 550894 549854 586338
rect 549234 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 549854 550894
rect 549234 550574 549854 550658
rect 549234 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 549854 550574
rect 549234 514894 549854 550338
rect 549234 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 549854 514894
rect 549234 514574 549854 514658
rect 549234 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 549854 514574
rect 549234 478894 549854 514338
rect 549234 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 549854 478894
rect 549234 478574 549854 478658
rect 549234 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 549854 478574
rect 549234 442894 549854 478338
rect 549234 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 549854 442894
rect 549234 442574 549854 442658
rect 549234 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 549854 442574
rect 549234 406894 549854 442338
rect 549234 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 549854 406894
rect 549234 406574 549854 406658
rect 549234 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 549854 406574
rect 549234 370894 549854 406338
rect 549234 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 549854 370894
rect 549234 370574 549854 370658
rect 549234 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 549854 370574
rect 549234 334894 549854 370338
rect 549234 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 549854 334894
rect 549234 334574 549854 334658
rect 549234 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 549854 334574
rect 549234 298894 549854 334338
rect 549234 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 549854 298894
rect 549234 298574 549854 298658
rect 549234 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 549854 298574
rect 549234 262894 549854 298338
rect 549234 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 549854 262894
rect 549234 262574 549854 262658
rect 549234 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 549854 262574
rect 549234 226894 549854 262338
rect 549234 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 549854 226894
rect 549234 226574 549854 226658
rect 549234 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 549854 226574
rect 549234 190894 549854 226338
rect 549234 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 549854 190894
rect 549234 190574 549854 190658
rect 549234 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 549854 190574
rect 549234 154894 549854 190338
rect 549234 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 549854 154894
rect 549234 154574 549854 154658
rect 549234 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 549854 154574
rect 549234 118894 549854 154338
rect 549234 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 549854 118894
rect 549234 118574 549854 118658
rect 549234 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 549854 118574
rect 549234 82894 549854 118338
rect 549234 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 549854 82894
rect 549234 82574 549854 82658
rect 549234 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 549854 82574
rect 549234 46894 549854 82338
rect 549234 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 549854 46894
rect 549234 46574 549854 46658
rect 549234 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 549854 46574
rect 549234 10894 549854 46338
rect 549234 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 549854 10894
rect 549234 10574 549854 10658
rect 549234 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 549854 10574
rect 549234 -4186 549854 10338
rect 549234 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 549854 -4186
rect 549234 -4506 549854 -4422
rect 549234 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 549854 -4506
rect 549234 -5734 549854 -4742
rect 552954 698614 553574 710042
rect 570954 711558 571574 711590
rect 570954 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 571574 711558
rect 570954 711238 571574 711322
rect 570954 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 571574 711238
rect 567234 709638 567854 709670
rect 567234 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 567854 709638
rect 567234 709318 567854 709402
rect 567234 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 567854 709318
rect 563514 707718 564134 707750
rect 563514 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 564134 707718
rect 563514 707398 564134 707482
rect 563514 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 564134 707398
rect 552954 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 553574 698614
rect 552954 698294 553574 698378
rect 552954 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 553574 698294
rect 552954 662614 553574 698058
rect 552954 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 553574 662614
rect 552954 662294 553574 662378
rect 552954 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 553574 662294
rect 552954 626614 553574 662058
rect 552954 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 553574 626614
rect 552954 626294 553574 626378
rect 552954 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 553574 626294
rect 552954 590614 553574 626058
rect 552954 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 553574 590614
rect 552954 590294 553574 590378
rect 552954 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 553574 590294
rect 552954 554614 553574 590058
rect 552954 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 553574 554614
rect 552954 554294 553574 554378
rect 552954 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 553574 554294
rect 552954 518614 553574 554058
rect 552954 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 553574 518614
rect 552954 518294 553574 518378
rect 552954 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 553574 518294
rect 552954 482614 553574 518058
rect 552954 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 553574 482614
rect 552954 482294 553574 482378
rect 552954 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 553574 482294
rect 552954 446614 553574 482058
rect 552954 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 553574 446614
rect 552954 446294 553574 446378
rect 552954 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 553574 446294
rect 552954 410614 553574 446058
rect 552954 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 553574 410614
rect 552954 410294 553574 410378
rect 552954 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 553574 410294
rect 552954 374614 553574 410058
rect 552954 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 553574 374614
rect 552954 374294 553574 374378
rect 552954 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 553574 374294
rect 552954 338614 553574 374058
rect 552954 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 553574 338614
rect 552954 338294 553574 338378
rect 552954 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 553574 338294
rect 552954 302614 553574 338058
rect 552954 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 553574 302614
rect 552954 302294 553574 302378
rect 552954 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 553574 302294
rect 552954 266614 553574 302058
rect 552954 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 553574 266614
rect 552954 266294 553574 266378
rect 552954 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 553574 266294
rect 552954 230614 553574 266058
rect 552954 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 553574 230614
rect 552954 230294 553574 230378
rect 552954 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 553574 230294
rect 552954 194614 553574 230058
rect 552954 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 553574 194614
rect 552954 194294 553574 194378
rect 552954 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 553574 194294
rect 552954 158614 553574 194058
rect 552954 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 553574 158614
rect 552954 158294 553574 158378
rect 552954 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 553574 158294
rect 552954 122614 553574 158058
rect 552954 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 553574 122614
rect 552954 122294 553574 122378
rect 552954 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 553574 122294
rect 552954 86614 553574 122058
rect 552954 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 553574 86614
rect 552954 86294 553574 86378
rect 552954 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 553574 86294
rect 552954 50614 553574 86058
rect 552954 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 553574 50614
rect 552954 50294 553574 50378
rect 552954 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 553574 50294
rect 552954 14614 553574 50058
rect 552954 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 553574 14614
rect 552954 14294 553574 14378
rect 552954 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 553574 14294
rect 534954 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 535574 -7066
rect 534954 -7386 535574 -7302
rect 534954 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 535574 -7386
rect 534954 -7654 535574 -7622
rect 552954 -6106 553574 14058
rect 559794 705798 560414 705830
rect 559794 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 560414 705798
rect 559794 705478 560414 705562
rect 559794 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 560414 705478
rect 559794 669454 560414 705242
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -1306 560414 20898
rect 559794 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 560414 -1306
rect 559794 -1626 560414 -1542
rect 559794 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 560414 -1626
rect 559794 -1894 560414 -1862
rect 563514 673174 564134 707162
rect 563514 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 564134 673174
rect 563514 672854 564134 672938
rect 563514 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 564134 672854
rect 563514 637174 564134 672618
rect 563514 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 564134 637174
rect 563514 636854 564134 636938
rect 563514 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 564134 636854
rect 563514 601174 564134 636618
rect 563514 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 564134 601174
rect 563514 600854 564134 600938
rect 563514 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 564134 600854
rect 563514 565174 564134 600618
rect 563514 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 564134 565174
rect 563514 564854 564134 564938
rect 563514 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 564134 564854
rect 563514 529174 564134 564618
rect 563514 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 564134 529174
rect 563514 528854 564134 528938
rect 563514 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 564134 528854
rect 563514 493174 564134 528618
rect 563514 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 564134 493174
rect 563514 492854 564134 492938
rect 563514 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 564134 492854
rect 563514 457174 564134 492618
rect 563514 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 564134 457174
rect 563514 456854 564134 456938
rect 563514 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 564134 456854
rect 563514 421174 564134 456618
rect 563514 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 564134 421174
rect 563514 420854 564134 420938
rect 563514 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 564134 420854
rect 563514 385174 564134 420618
rect 563514 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 564134 385174
rect 563514 384854 564134 384938
rect 563514 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 564134 384854
rect 563514 349174 564134 384618
rect 563514 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 564134 349174
rect 563514 348854 564134 348938
rect 563514 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 564134 348854
rect 563514 313174 564134 348618
rect 563514 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 564134 313174
rect 563514 312854 564134 312938
rect 563514 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 564134 312854
rect 563514 277174 564134 312618
rect 563514 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 564134 277174
rect 563514 276854 564134 276938
rect 563514 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 564134 276854
rect 563514 241174 564134 276618
rect 563514 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 564134 241174
rect 563514 240854 564134 240938
rect 563514 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 564134 240854
rect 563514 205174 564134 240618
rect 563514 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 564134 205174
rect 563514 204854 564134 204938
rect 563514 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 564134 204854
rect 563514 169174 564134 204618
rect 563514 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 564134 169174
rect 563514 168854 564134 168938
rect 563514 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 564134 168854
rect 563514 133174 564134 168618
rect 563514 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 564134 133174
rect 563514 132854 564134 132938
rect 563514 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 564134 132854
rect 563514 97174 564134 132618
rect 563514 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 564134 97174
rect 563514 96854 564134 96938
rect 563514 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 564134 96854
rect 563514 61174 564134 96618
rect 563514 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 564134 61174
rect 563514 60854 564134 60938
rect 563514 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 564134 60854
rect 563514 25174 564134 60618
rect 563514 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 564134 25174
rect 563514 24854 564134 24938
rect 563514 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 564134 24854
rect 563514 -3226 564134 24618
rect 563514 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 564134 -3226
rect 563514 -3546 564134 -3462
rect 563514 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 564134 -3546
rect 563514 -3814 564134 -3782
rect 567234 676894 567854 709082
rect 567234 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 567854 676894
rect 567234 676574 567854 676658
rect 567234 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 567854 676574
rect 567234 640894 567854 676338
rect 567234 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 567854 640894
rect 567234 640574 567854 640658
rect 567234 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 567854 640574
rect 567234 604894 567854 640338
rect 567234 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 567854 604894
rect 567234 604574 567854 604658
rect 567234 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 567854 604574
rect 567234 568894 567854 604338
rect 567234 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 567854 568894
rect 567234 568574 567854 568658
rect 567234 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 567854 568574
rect 567234 532894 567854 568338
rect 567234 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 567854 532894
rect 567234 532574 567854 532658
rect 567234 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 567854 532574
rect 567234 496894 567854 532338
rect 567234 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 567854 496894
rect 567234 496574 567854 496658
rect 567234 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 567854 496574
rect 567234 460894 567854 496338
rect 567234 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 567854 460894
rect 567234 460574 567854 460658
rect 567234 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 567854 460574
rect 567234 424894 567854 460338
rect 567234 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 567854 424894
rect 567234 424574 567854 424658
rect 567234 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 567854 424574
rect 567234 388894 567854 424338
rect 567234 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 567854 388894
rect 567234 388574 567854 388658
rect 567234 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 567854 388574
rect 567234 352894 567854 388338
rect 567234 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 567854 352894
rect 567234 352574 567854 352658
rect 567234 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 567854 352574
rect 567234 316894 567854 352338
rect 567234 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 567854 316894
rect 567234 316574 567854 316658
rect 567234 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 567854 316574
rect 567234 280894 567854 316338
rect 567234 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 567854 280894
rect 567234 280574 567854 280658
rect 567234 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 567854 280574
rect 567234 244894 567854 280338
rect 567234 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 567854 244894
rect 567234 244574 567854 244658
rect 567234 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 567854 244574
rect 567234 208894 567854 244338
rect 567234 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 567854 208894
rect 567234 208574 567854 208658
rect 567234 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 567854 208574
rect 567234 172894 567854 208338
rect 567234 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 567854 172894
rect 567234 172574 567854 172658
rect 567234 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 567854 172574
rect 567234 136894 567854 172338
rect 567234 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 567854 136894
rect 567234 136574 567854 136658
rect 567234 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 567854 136574
rect 567234 100894 567854 136338
rect 567234 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 567854 100894
rect 567234 100574 567854 100658
rect 567234 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 567854 100574
rect 567234 64894 567854 100338
rect 567234 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 567854 64894
rect 567234 64574 567854 64658
rect 567234 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 567854 64574
rect 567234 28894 567854 64338
rect 567234 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 567854 28894
rect 567234 28574 567854 28658
rect 567234 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 567854 28574
rect 567234 -5146 567854 28338
rect 567234 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 567854 -5146
rect 567234 -5466 567854 -5382
rect 567234 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 567854 -5466
rect 567234 -5734 567854 -5702
rect 570954 680614 571574 711002
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 581514 706758 582134 707750
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 581514 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 582134 706758
rect 581514 706438 582134 706522
rect 581514 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 582134 706438
rect 570954 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 571574 680614
rect 570954 680294 571574 680378
rect 570954 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 571574 680294
rect 570954 644614 571574 680058
rect 570954 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 571574 644614
rect 570954 644294 571574 644378
rect 570954 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 571574 644294
rect 570954 608614 571574 644058
rect 570954 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 571574 608614
rect 570954 608294 571574 608378
rect 570954 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 571574 608294
rect 570954 572614 571574 608058
rect 570954 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 571574 572614
rect 570954 572294 571574 572378
rect 570954 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 571574 572294
rect 570954 536614 571574 572058
rect 570954 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 571574 536614
rect 570954 536294 571574 536378
rect 570954 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 571574 536294
rect 570954 500614 571574 536058
rect 570954 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 571574 500614
rect 570954 500294 571574 500378
rect 570954 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 571574 500294
rect 570954 464614 571574 500058
rect 570954 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 571574 464614
rect 570954 464294 571574 464378
rect 570954 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 571574 464294
rect 570954 428614 571574 464058
rect 570954 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 571574 428614
rect 570954 428294 571574 428378
rect 570954 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 571574 428294
rect 570954 392614 571574 428058
rect 570954 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 571574 392614
rect 570954 392294 571574 392378
rect 570954 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 571574 392294
rect 570954 356614 571574 392058
rect 570954 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 571574 356614
rect 570954 356294 571574 356378
rect 570954 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 571574 356294
rect 570954 320614 571574 356058
rect 570954 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 571574 320614
rect 570954 320294 571574 320378
rect 570954 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 571574 320294
rect 570954 284614 571574 320058
rect 570954 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 571574 284614
rect 570954 284294 571574 284378
rect 570954 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 571574 284294
rect 570954 248614 571574 284058
rect 570954 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 571574 248614
rect 570954 248294 571574 248378
rect 570954 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 571574 248294
rect 570954 212614 571574 248058
rect 570954 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 571574 212614
rect 570954 212294 571574 212378
rect 570954 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 571574 212294
rect 570954 176614 571574 212058
rect 570954 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 571574 176614
rect 570954 176294 571574 176378
rect 570954 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 571574 176294
rect 570954 140614 571574 176058
rect 570954 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 571574 140614
rect 570954 140294 571574 140378
rect 570954 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 571574 140294
rect 570954 104614 571574 140058
rect 570954 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 571574 104614
rect 570954 104294 571574 104378
rect 570954 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 571574 104294
rect 570954 68614 571574 104058
rect 570954 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 571574 68614
rect 570954 68294 571574 68378
rect 570954 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 571574 68294
rect 570954 32614 571574 68058
rect 570954 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 571574 32614
rect 570954 32294 571574 32378
rect 570954 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 571574 32294
rect 552954 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 553574 -6106
rect 552954 -6426 553574 -6342
rect 552954 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 553574 -6426
rect 552954 -7654 553574 -6662
rect 570954 -7066 571574 32058
rect 577794 704838 578414 705830
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 580211 697236 580277 697237
rect 580211 697172 580212 697236
rect 580276 697172 580277 697236
rect 580211 697171 580277 697172
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 580214 179077 580274 697171
rect 581514 691174 582134 706202
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 580395 683908 580461 683909
rect 580395 683844 580396 683908
rect 580460 683844 580461 683908
rect 580395 683843 580461 683844
rect 580211 179076 580277 179077
rect 580211 179012 580212 179076
rect 580276 179012 580277 179076
rect 580211 179011 580277 179012
rect 580398 178669 580458 683843
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 580579 630868 580645 630869
rect 580579 630804 580580 630868
rect 580644 630804 580645 630868
rect 580579 630803 580645 630804
rect 580582 179485 580642 630803
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 580579 179484 580645 179485
rect 580579 179420 580580 179484
rect 580644 179420 580645 179484
rect 580579 179419 580645 179420
rect 580395 178668 580461 178669
rect 580395 178604 580396 178668
rect 580460 178604 580461 178668
rect 580395 178603 580461 178604
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -1894 578414 -902
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -2266 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 669454 586890 705242
rect 586270 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect 586270 669134 586890 669218
rect 586270 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect 586270 633454 586890 668898
rect 586270 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect 586270 633134 586890 633218
rect 586270 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect 586270 597454 586890 632898
rect 586270 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect 586270 597134 586890 597218
rect 586270 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect 586270 561454 586890 596898
rect 586270 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect 586270 561134 586890 561218
rect 586270 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect 586270 525454 586890 560898
rect 586270 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect 586270 525134 586890 525218
rect 586270 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect 586270 489454 586890 524898
rect 586270 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect 586270 489134 586890 489218
rect 586270 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect 586270 453454 586890 488898
rect 586270 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect 586270 453134 586890 453218
rect 586270 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect 586270 417454 586890 452898
rect 586270 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect 586270 417134 586890 417218
rect 586270 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect 586270 381454 586890 416898
rect 586270 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect 586270 381134 586890 381218
rect 586270 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect 586270 345454 586890 380898
rect 586270 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect 586270 345134 586890 345218
rect 586270 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect 586270 309454 586890 344898
rect 586270 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect 586270 309134 586890 309218
rect 586270 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect 586270 273454 586890 308898
rect 586270 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect 586270 273134 586890 273218
rect 586270 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect 586270 237454 586890 272898
rect 586270 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect 586270 237134 586890 237218
rect 586270 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect 586270 201454 586890 236898
rect 586270 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect 586270 201134 586890 201218
rect 586270 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect 586270 165454 586890 200898
rect 586270 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect 586270 165134 586890 165218
rect 586270 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect 586270 129454 586890 164898
rect 586270 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect 586270 129134 586890 129218
rect 586270 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect 586270 93454 586890 128898
rect 586270 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect 586270 93134 586890 93218
rect 586270 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect 586270 57454 586890 92898
rect 586270 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect 586270 57134 586890 57218
rect 586270 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect 586270 21454 586890 56898
rect 586270 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect 586270 21134 586890 21218
rect 586270 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect 586270 -1306 586890 20898
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 691174 587850 706202
rect 587230 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 587850 691174
rect 587230 690854 587850 690938
rect 587230 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 587850 690854
rect 587230 655174 587850 690618
rect 587230 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 587850 655174
rect 587230 654854 587850 654938
rect 587230 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 587850 654854
rect 587230 619174 587850 654618
rect 587230 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 587850 619174
rect 587230 618854 587850 618938
rect 587230 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 587850 618854
rect 587230 583174 587850 618618
rect 587230 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 587850 583174
rect 587230 582854 587850 582938
rect 587230 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 587850 582854
rect 587230 547174 587850 582618
rect 587230 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 587850 547174
rect 587230 546854 587850 546938
rect 587230 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 587850 546854
rect 587230 511174 587850 546618
rect 587230 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 587850 511174
rect 587230 510854 587850 510938
rect 587230 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 587850 510854
rect 587230 475174 587850 510618
rect 587230 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 587850 475174
rect 587230 474854 587850 474938
rect 587230 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 587850 474854
rect 587230 439174 587850 474618
rect 587230 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 587850 439174
rect 587230 438854 587850 438938
rect 587230 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 587850 438854
rect 587230 403174 587850 438618
rect 587230 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 587850 403174
rect 587230 402854 587850 402938
rect 587230 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 587850 402854
rect 587230 367174 587850 402618
rect 587230 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 587850 367174
rect 587230 366854 587850 366938
rect 587230 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 587850 366854
rect 587230 331174 587850 366618
rect 587230 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 587850 331174
rect 587230 330854 587850 330938
rect 587230 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 587850 330854
rect 587230 295174 587850 330618
rect 587230 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 587850 295174
rect 587230 294854 587850 294938
rect 587230 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 587850 294854
rect 587230 259174 587850 294618
rect 587230 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 587850 259174
rect 587230 258854 587850 258938
rect 587230 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 587850 258854
rect 587230 223174 587850 258618
rect 587230 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 587850 223174
rect 587230 222854 587850 222938
rect 587230 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 587850 222854
rect 587230 187174 587850 222618
rect 587230 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 587850 187174
rect 587230 186854 587850 186938
rect 587230 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 587850 186854
rect 587230 151174 587850 186618
rect 587230 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 587850 151174
rect 587230 150854 587850 150938
rect 587230 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 587850 150854
rect 587230 115174 587850 150618
rect 587230 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 587850 115174
rect 587230 114854 587850 114938
rect 587230 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 587850 114854
rect 587230 79174 587850 114618
rect 587230 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 587850 79174
rect 587230 78854 587850 78938
rect 587230 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 587850 78854
rect 587230 43174 587850 78618
rect 587230 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 587850 43174
rect 587230 42854 587850 42938
rect 587230 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 587850 42854
rect 587230 7174 587850 42618
rect 587230 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 587850 7174
rect 587230 6854 587850 6938
rect 587230 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 587850 6854
rect 581514 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 582134 -2266
rect 581514 -2586 582134 -2502
rect 581514 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 582134 -2586
rect 581514 -3814 582134 -2822
rect 587230 -2266 587850 6618
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 673174 588810 707162
rect 588190 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect 588190 672854 588810 672938
rect 588190 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect 588190 637174 588810 672618
rect 588190 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect 588190 636854 588810 636938
rect 588190 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect 588190 601174 588810 636618
rect 588190 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect 588190 600854 588810 600938
rect 588190 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect 588190 565174 588810 600618
rect 588190 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect 588190 564854 588810 564938
rect 588190 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect 588190 529174 588810 564618
rect 588190 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect 588190 528854 588810 528938
rect 588190 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect 588190 493174 588810 528618
rect 588190 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect 588190 492854 588810 492938
rect 588190 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect 588190 457174 588810 492618
rect 588190 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect 588190 456854 588810 456938
rect 588190 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect 588190 421174 588810 456618
rect 588190 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect 588190 420854 588810 420938
rect 588190 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect 588190 385174 588810 420618
rect 588190 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect 588190 384854 588810 384938
rect 588190 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect 588190 349174 588810 384618
rect 588190 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect 588190 348854 588810 348938
rect 588190 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect 588190 313174 588810 348618
rect 588190 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect 588190 312854 588810 312938
rect 588190 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect 588190 277174 588810 312618
rect 588190 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect 588190 276854 588810 276938
rect 588190 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect 588190 241174 588810 276618
rect 588190 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect 588190 240854 588810 240938
rect 588190 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect 588190 205174 588810 240618
rect 588190 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect 588190 204854 588810 204938
rect 588190 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect 588190 169174 588810 204618
rect 588190 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect 588190 168854 588810 168938
rect 588190 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect 588190 133174 588810 168618
rect 588190 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect 588190 132854 588810 132938
rect 588190 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect 588190 97174 588810 132618
rect 588190 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect 588190 96854 588810 96938
rect 588190 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect 588190 61174 588810 96618
rect 588190 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect 588190 60854 588810 60938
rect 588190 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect 588190 25174 588810 60618
rect 588190 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect 588190 24854 588810 24938
rect 588190 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect 588190 -3226 588810 24618
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 694894 589770 708122
rect 589150 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 589770 694894
rect 589150 694574 589770 694658
rect 589150 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 589770 694574
rect 589150 658894 589770 694338
rect 589150 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 589770 658894
rect 589150 658574 589770 658658
rect 589150 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 589770 658574
rect 589150 622894 589770 658338
rect 589150 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 589770 622894
rect 589150 622574 589770 622658
rect 589150 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 589770 622574
rect 589150 586894 589770 622338
rect 589150 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 589770 586894
rect 589150 586574 589770 586658
rect 589150 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 589770 586574
rect 589150 550894 589770 586338
rect 589150 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 589770 550894
rect 589150 550574 589770 550658
rect 589150 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 589770 550574
rect 589150 514894 589770 550338
rect 589150 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 589770 514894
rect 589150 514574 589770 514658
rect 589150 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 589770 514574
rect 589150 478894 589770 514338
rect 589150 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 589770 478894
rect 589150 478574 589770 478658
rect 589150 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 589770 478574
rect 589150 442894 589770 478338
rect 589150 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 589770 442894
rect 589150 442574 589770 442658
rect 589150 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 589770 442574
rect 589150 406894 589770 442338
rect 589150 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 589770 406894
rect 589150 406574 589770 406658
rect 589150 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 589770 406574
rect 589150 370894 589770 406338
rect 589150 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 589770 370894
rect 589150 370574 589770 370658
rect 589150 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 589770 370574
rect 589150 334894 589770 370338
rect 589150 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 589770 334894
rect 589150 334574 589770 334658
rect 589150 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 589770 334574
rect 589150 298894 589770 334338
rect 589150 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 589770 298894
rect 589150 298574 589770 298658
rect 589150 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 589770 298574
rect 589150 262894 589770 298338
rect 589150 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 589770 262894
rect 589150 262574 589770 262658
rect 589150 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 589770 262574
rect 589150 226894 589770 262338
rect 589150 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 589770 226894
rect 589150 226574 589770 226658
rect 589150 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 589770 226574
rect 589150 190894 589770 226338
rect 589150 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 589770 190894
rect 589150 190574 589770 190658
rect 589150 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 589770 190574
rect 589150 154894 589770 190338
rect 589150 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 589770 154894
rect 589150 154574 589770 154658
rect 589150 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 589770 154574
rect 589150 118894 589770 154338
rect 589150 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 589770 118894
rect 589150 118574 589770 118658
rect 589150 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 589770 118574
rect 589150 82894 589770 118338
rect 589150 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 589770 82894
rect 589150 82574 589770 82658
rect 589150 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 589770 82574
rect 589150 46894 589770 82338
rect 589150 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 589770 46894
rect 589150 46574 589770 46658
rect 589150 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 589770 46574
rect 589150 10894 589770 46338
rect 589150 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 589770 10894
rect 589150 10574 589770 10658
rect 589150 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 589770 10574
rect 589150 -4186 589770 10338
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 676894 590730 709082
rect 590110 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect 590110 676574 590730 676658
rect 590110 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect 590110 640894 590730 676338
rect 590110 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect 590110 640574 590730 640658
rect 590110 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect 590110 604894 590730 640338
rect 590110 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect 590110 604574 590730 604658
rect 590110 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect 590110 568894 590730 604338
rect 590110 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect 590110 568574 590730 568658
rect 590110 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect 590110 532894 590730 568338
rect 590110 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect 590110 532574 590730 532658
rect 590110 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect 590110 496894 590730 532338
rect 590110 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect 590110 496574 590730 496658
rect 590110 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect 590110 460894 590730 496338
rect 590110 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect 590110 460574 590730 460658
rect 590110 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect 590110 424894 590730 460338
rect 590110 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect 590110 424574 590730 424658
rect 590110 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect 590110 388894 590730 424338
rect 590110 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect 590110 388574 590730 388658
rect 590110 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect 590110 352894 590730 388338
rect 590110 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect 590110 352574 590730 352658
rect 590110 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect 590110 316894 590730 352338
rect 590110 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect 590110 316574 590730 316658
rect 590110 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect 590110 280894 590730 316338
rect 590110 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect 590110 280574 590730 280658
rect 590110 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect 590110 244894 590730 280338
rect 590110 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect 590110 244574 590730 244658
rect 590110 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect 590110 208894 590730 244338
rect 590110 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect 590110 208574 590730 208658
rect 590110 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect 590110 172894 590730 208338
rect 590110 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect 590110 172574 590730 172658
rect 590110 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect 590110 136894 590730 172338
rect 590110 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect 590110 136574 590730 136658
rect 590110 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect 590110 100894 590730 136338
rect 590110 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect 590110 100574 590730 100658
rect 590110 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect 590110 64894 590730 100338
rect 590110 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect 590110 64574 590730 64658
rect 590110 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect 590110 28894 590730 64338
rect 590110 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect 590110 28574 590730 28658
rect 590110 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect 590110 -5146 590730 28338
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 698614 591690 710042
rect 591070 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 591690 698614
rect 591070 698294 591690 698378
rect 591070 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 591690 698294
rect 591070 662614 591690 698058
rect 591070 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 591690 662614
rect 591070 662294 591690 662378
rect 591070 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 591690 662294
rect 591070 626614 591690 662058
rect 591070 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 591690 626614
rect 591070 626294 591690 626378
rect 591070 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 591690 626294
rect 591070 590614 591690 626058
rect 591070 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 591690 590614
rect 591070 590294 591690 590378
rect 591070 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 591690 590294
rect 591070 554614 591690 590058
rect 591070 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 591690 554614
rect 591070 554294 591690 554378
rect 591070 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 591690 554294
rect 591070 518614 591690 554058
rect 591070 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 591690 518614
rect 591070 518294 591690 518378
rect 591070 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 591690 518294
rect 591070 482614 591690 518058
rect 591070 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 591690 482614
rect 591070 482294 591690 482378
rect 591070 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 591690 482294
rect 591070 446614 591690 482058
rect 591070 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 591690 446614
rect 591070 446294 591690 446378
rect 591070 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 591690 446294
rect 591070 410614 591690 446058
rect 591070 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 591690 410614
rect 591070 410294 591690 410378
rect 591070 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 591690 410294
rect 591070 374614 591690 410058
rect 591070 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 591690 374614
rect 591070 374294 591690 374378
rect 591070 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 591690 374294
rect 591070 338614 591690 374058
rect 591070 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 591690 338614
rect 591070 338294 591690 338378
rect 591070 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 591690 338294
rect 591070 302614 591690 338058
rect 591070 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 591690 302614
rect 591070 302294 591690 302378
rect 591070 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 591690 302294
rect 591070 266614 591690 302058
rect 591070 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 591690 266614
rect 591070 266294 591690 266378
rect 591070 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 591690 266294
rect 591070 230614 591690 266058
rect 591070 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 591690 230614
rect 591070 230294 591690 230378
rect 591070 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 591690 230294
rect 591070 194614 591690 230058
rect 591070 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 591690 194614
rect 591070 194294 591690 194378
rect 591070 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 591690 194294
rect 591070 158614 591690 194058
rect 591070 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 591690 158614
rect 591070 158294 591690 158378
rect 591070 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 591690 158294
rect 591070 122614 591690 158058
rect 591070 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 591690 122614
rect 591070 122294 591690 122378
rect 591070 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 591690 122294
rect 591070 86614 591690 122058
rect 591070 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 591690 86614
rect 591070 86294 591690 86378
rect 591070 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 591690 86294
rect 591070 50614 591690 86058
rect 591070 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 591690 50614
rect 591070 50294 591690 50378
rect 591070 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 591690 50294
rect 591070 14614 591690 50058
rect 591070 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 591690 14614
rect 591070 14294 591690 14378
rect 591070 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 591690 14294
rect 591070 -6106 591690 14058
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 680614 592650 711002
rect 592030 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect 592030 680294 592650 680378
rect 592030 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect 592030 644614 592650 680058
rect 592030 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect 592030 644294 592650 644378
rect 592030 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect 592030 608614 592650 644058
rect 592030 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect 592030 608294 592650 608378
rect 592030 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect 592030 572614 592650 608058
rect 592030 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect 592030 572294 592650 572378
rect 592030 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect 592030 536614 592650 572058
rect 592030 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect 592030 536294 592650 536378
rect 592030 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect 592030 500614 592650 536058
rect 592030 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect 592030 500294 592650 500378
rect 592030 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect 592030 464614 592650 500058
rect 592030 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect 592030 464294 592650 464378
rect 592030 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect 592030 428614 592650 464058
rect 592030 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect 592030 428294 592650 428378
rect 592030 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect 592030 392614 592650 428058
rect 592030 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect 592030 392294 592650 392378
rect 592030 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect 592030 356614 592650 392058
rect 592030 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect 592030 356294 592650 356378
rect 592030 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect 592030 320614 592650 356058
rect 592030 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect 592030 320294 592650 320378
rect 592030 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect 592030 284614 592650 320058
rect 592030 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect 592030 284294 592650 284378
rect 592030 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect 592030 248614 592650 284058
rect 592030 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect 592030 248294 592650 248378
rect 592030 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect 592030 212614 592650 248058
rect 592030 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect 592030 212294 592650 212378
rect 592030 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect 592030 176614 592650 212058
rect 592030 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect 592030 176294 592650 176378
rect 592030 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect 592030 140614 592650 176058
rect 592030 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect 592030 140294 592650 140378
rect 592030 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect 592030 104614 592650 140058
rect 592030 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect 592030 104294 592650 104378
rect 592030 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect 592030 68614 592650 104058
rect 592030 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect 592030 68294 592650 68378
rect 592030 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect 592030 32614 592650 68058
rect 592030 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect 592030 32294 592650 32378
rect 592030 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect 570954 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 571574 -7066
rect 570954 -7386 571574 -7302
rect 570954 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 571574 -7386
rect 570954 -7654 571574 -7622
rect 592030 -7066 592650 32058
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 680378 -8458 680614
rect -8374 680378 -8138 680614
rect -8694 680058 -8458 680294
rect -8374 680058 -8138 680294
rect -8694 644378 -8458 644614
rect -8374 644378 -8138 644614
rect -8694 644058 -8458 644294
rect -8374 644058 -8138 644294
rect -8694 608378 -8458 608614
rect -8374 608378 -8138 608614
rect -8694 608058 -8458 608294
rect -8374 608058 -8138 608294
rect -8694 572378 -8458 572614
rect -8374 572378 -8138 572614
rect -8694 572058 -8458 572294
rect -8374 572058 -8138 572294
rect -8694 536378 -8458 536614
rect -8374 536378 -8138 536614
rect -8694 536058 -8458 536294
rect -8374 536058 -8138 536294
rect -8694 500378 -8458 500614
rect -8374 500378 -8138 500614
rect -8694 500058 -8458 500294
rect -8374 500058 -8138 500294
rect -8694 464378 -8458 464614
rect -8374 464378 -8138 464614
rect -8694 464058 -8458 464294
rect -8374 464058 -8138 464294
rect -8694 428378 -8458 428614
rect -8374 428378 -8138 428614
rect -8694 428058 -8458 428294
rect -8374 428058 -8138 428294
rect -8694 392378 -8458 392614
rect -8374 392378 -8138 392614
rect -8694 392058 -8458 392294
rect -8374 392058 -8138 392294
rect -8694 356378 -8458 356614
rect -8374 356378 -8138 356614
rect -8694 356058 -8458 356294
rect -8374 356058 -8138 356294
rect -8694 320378 -8458 320614
rect -8374 320378 -8138 320614
rect -8694 320058 -8458 320294
rect -8374 320058 -8138 320294
rect -8694 284378 -8458 284614
rect -8374 284378 -8138 284614
rect -8694 284058 -8458 284294
rect -8374 284058 -8138 284294
rect -8694 248378 -8458 248614
rect -8374 248378 -8138 248614
rect -8694 248058 -8458 248294
rect -8374 248058 -8138 248294
rect -8694 212378 -8458 212614
rect -8374 212378 -8138 212614
rect -8694 212058 -8458 212294
rect -8374 212058 -8138 212294
rect -8694 176378 -8458 176614
rect -8374 176378 -8138 176614
rect -8694 176058 -8458 176294
rect -8374 176058 -8138 176294
rect -8694 140378 -8458 140614
rect -8374 140378 -8138 140614
rect -8694 140058 -8458 140294
rect -8374 140058 -8138 140294
rect -8694 104378 -8458 104614
rect -8374 104378 -8138 104614
rect -8694 104058 -8458 104294
rect -8374 104058 -8138 104294
rect -8694 68378 -8458 68614
rect -8374 68378 -8138 68614
rect -8694 68058 -8458 68294
rect -8374 68058 -8138 68294
rect -8694 32378 -8458 32614
rect -8374 32378 -8138 32614
rect -8694 32058 -8458 32294
rect -8374 32058 -8138 32294
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect 12986 710362 13222 710598
rect 13306 710362 13542 710598
rect 12986 710042 13222 710278
rect 13306 710042 13542 710278
rect -7734 698378 -7498 698614
rect -7414 698378 -7178 698614
rect -7734 698058 -7498 698294
rect -7414 698058 -7178 698294
rect -7734 662378 -7498 662614
rect -7414 662378 -7178 662614
rect -7734 662058 -7498 662294
rect -7414 662058 -7178 662294
rect -7734 626378 -7498 626614
rect -7414 626378 -7178 626614
rect -7734 626058 -7498 626294
rect -7414 626058 -7178 626294
rect -7734 590378 -7498 590614
rect -7414 590378 -7178 590614
rect -7734 590058 -7498 590294
rect -7414 590058 -7178 590294
rect -7734 554378 -7498 554614
rect -7414 554378 -7178 554614
rect -7734 554058 -7498 554294
rect -7414 554058 -7178 554294
rect -7734 518378 -7498 518614
rect -7414 518378 -7178 518614
rect -7734 518058 -7498 518294
rect -7414 518058 -7178 518294
rect -7734 482378 -7498 482614
rect -7414 482378 -7178 482614
rect -7734 482058 -7498 482294
rect -7414 482058 -7178 482294
rect -7734 446378 -7498 446614
rect -7414 446378 -7178 446614
rect -7734 446058 -7498 446294
rect -7414 446058 -7178 446294
rect -7734 410378 -7498 410614
rect -7414 410378 -7178 410614
rect -7734 410058 -7498 410294
rect -7414 410058 -7178 410294
rect -7734 374378 -7498 374614
rect -7414 374378 -7178 374614
rect -7734 374058 -7498 374294
rect -7414 374058 -7178 374294
rect -7734 338378 -7498 338614
rect -7414 338378 -7178 338614
rect -7734 338058 -7498 338294
rect -7414 338058 -7178 338294
rect -7734 302378 -7498 302614
rect -7414 302378 -7178 302614
rect -7734 302058 -7498 302294
rect -7414 302058 -7178 302294
rect -7734 266378 -7498 266614
rect -7414 266378 -7178 266614
rect -7734 266058 -7498 266294
rect -7414 266058 -7178 266294
rect -7734 230378 -7498 230614
rect -7414 230378 -7178 230614
rect -7734 230058 -7498 230294
rect -7414 230058 -7178 230294
rect -7734 194378 -7498 194614
rect -7414 194378 -7178 194614
rect -7734 194058 -7498 194294
rect -7414 194058 -7178 194294
rect -7734 158378 -7498 158614
rect -7414 158378 -7178 158614
rect -7734 158058 -7498 158294
rect -7414 158058 -7178 158294
rect -7734 122378 -7498 122614
rect -7414 122378 -7178 122614
rect -7734 122058 -7498 122294
rect -7414 122058 -7178 122294
rect -7734 86378 -7498 86614
rect -7414 86378 -7178 86614
rect -7734 86058 -7498 86294
rect -7414 86058 -7178 86294
rect -7734 50378 -7498 50614
rect -7414 50378 -7178 50614
rect -7734 50058 -7498 50294
rect -7414 50058 -7178 50294
rect -7734 14378 -7498 14614
rect -7414 14378 -7178 14614
rect -7734 14058 -7498 14294
rect -7414 14058 -7178 14294
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 676658 -6538 676894
rect -6454 676658 -6218 676894
rect -6774 676338 -6538 676574
rect -6454 676338 -6218 676574
rect -6774 640658 -6538 640894
rect -6454 640658 -6218 640894
rect -6774 640338 -6538 640574
rect -6454 640338 -6218 640574
rect -6774 604658 -6538 604894
rect -6454 604658 -6218 604894
rect -6774 604338 -6538 604574
rect -6454 604338 -6218 604574
rect -6774 568658 -6538 568894
rect -6454 568658 -6218 568894
rect -6774 568338 -6538 568574
rect -6454 568338 -6218 568574
rect -6774 532658 -6538 532894
rect -6454 532658 -6218 532894
rect -6774 532338 -6538 532574
rect -6454 532338 -6218 532574
rect -6774 496658 -6538 496894
rect -6454 496658 -6218 496894
rect -6774 496338 -6538 496574
rect -6454 496338 -6218 496574
rect -6774 460658 -6538 460894
rect -6454 460658 -6218 460894
rect -6774 460338 -6538 460574
rect -6454 460338 -6218 460574
rect -6774 424658 -6538 424894
rect -6454 424658 -6218 424894
rect -6774 424338 -6538 424574
rect -6454 424338 -6218 424574
rect -6774 388658 -6538 388894
rect -6454 388658 -6218 388894
rect -6774 388338 -6538 388574
rect -6454 388338 -6218 388574
rect -6774 352658 -6538 352894
rect -6454 352658 -6218 352894
rect -6774 352338 -6538 352574
rect -6454 352338 -6218 352574
rect -6774 316658 -6538 316894
rect -6454 316658 -6218 316894
rect -6774 316338 -6538 316574
rect -6454 316338 -6218 316574
rect -6774 280658 -6538 280894
rect -6454 280658 -6218 280894
rect -6774 280338 -6538 280574
rect -6454 280338 -6218 280574
rect -6774 244658 -6538 244894
rect -6454 244658 -6218 244894
rect -6774 244338 -6538 244574
rect -6454 244338 -6218 244574
rect -6774 208658 -6538 208894
rect -6454 208658 -6218 208894
rect -6774 208338 -6538 208574
rect -6454 208338 -6218 208574
rect -6774 172658 -6538 172894
rect -6454 172658 -6218 172894
rect -6774 172338 -6538 172574
rect -6454 172338 -6218 172574
rect -6774 136658 -6538 136894
rect -6454 136658 -6218 136894
rect -6774 136338 -6538 136574
rect -6454 136338 -6218 136574
rect -6774 100658 -6538 100894
rect -6454 100658 -6218 100894
rect -6774 100338 -6538 100574
rect -6454 100338 -6218 100574
rect -6774 64658 -6538 64894
rect -6454 64658 -6218 64894
rect -6774 64338 -6538 64574
rect -6454 64338 -6218 64574
rect -6774 28658 -6538 28894
rect -6454 28658 -6218 28894
rect -6774 28338 -6538 28574
rect -6454 28338 -6218 28574
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect 9266 708442 9502 708678
rect 9586 708442 9822 708678
rect 9266 708122 9502 708358
rect 9586 708122 9822 708358
rect -5814 694658 -5578 694894
rect -5494 694658 -5258 694894
rect -5814 694338 -5578 694574
rect -5494 694338 -5258 694574
rect -5814 658658 -5578 658894
rect -5494 658658 -5258 658894
rect -5814 658338 -5578 658574
rect -5494 658338 -5258 658574
rect -5814 622658 -5578 622894
rect -5494 622658 -5258 622894
rect -5814 622338 -5578 622574
rect -5494 622338 -5258 622574
rect -5814 586658 -5578 586894
rect -5494 586658 -5258 586894
rect -5814 586338 -5578 586574
rect -5494 586338 -5258 586574
rect -5814 550658 -5578 550894
rect -5494 550658 -5258 550894
rect -5814 550338 -5578 550574
rect -5494 550338 -5258 550574
rect -5814 514658 -5578 514894
rect -5494 514658 -5258 514894
rect -5814 514338 -5578 514574
rect -5494 514338 -5258 514574
rect -5814 478658 -5578 478894
rect -5494 478658 -5258 478894
rect -5814 478338 -5578 478574
rect -5494 478338 -5258 478574
rect -5814 442658 -5578 442894
rect -5494 442658 -5258 442894
rect -5814 442338 -5578 442574
rect -5494 442338 -5258 442574
rect -5814 406658 -5578 406894
rect -5494 406658 -5258 406894
rect -5814 406338 -5578 406574
rect -5494 406338 -5258 406574
rect -5814 370658 -5578 370894
rect -5494 370658 -5258 370894
rect -5814 370338 -5578 370574
rect -5494 370338 -5258 370574
rect -5814 334658 -5578 334894
rect -5494 334658 -5258 334894
rect -5814 334338 -5578 334574
rect -5494 334338 -5258 334574
rect -5814 298658 -5578 298894
rect -5494 298658 -5258 298894
rect -5814 298338 -5578 298574
rect -5494 298338 -5258 298574
rect -5814 262658 -5578 262894
rect -5494 262658 -5258 262894
rect -5814 262338 -5578 262574
rect -5494 262338 -5258 262574
rect -5814 226658 -5578 226894
rect -5494 226658 -5258 226894
rect -5814 226338 -5578 226574
rect -5494 226338 -5258 226574
rect -5814 190658 -5578 190894
rect -5494 190658 -5258 190894
rect -5814 190338 -5578 190574
rect -5494 190338 -5258 190574
rect -5814 154658 -5578 154894
rect -5494 154658 -5258 154894
rect -5814 154338 -5578 154574
rect -5494 154338 -5258 154574
rect -5814 118658 -5578 118894
rect -5494 118658 -5258 118894
rect -5814 118338 -5578 118574
rect -5494 118338 -5258 118574
rect -5814 82658 -5578 82894
rect -5494 82658 -5258 82894
rect -5814 82338 -5578 82574
rect -5494 82338 -5258 82574
rect -5814 46658 -5578 46894
rect -5494 46658 -5258 46894
rect -5814 46338 -5578 46574
rect -5494 46338 -5258 46574
rect -5814 10658 -5578 10894
rect -5494 10658 -5258 10894
rect -5814 10338 -5578 10574
rect -5494 10338 -5258 10574
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 672938 -4618 673174
rect -4534 672938 -4298 673174
rect -4854 672618 -4618 672854
rect -4534 672618 -4298 672854
rect -4854 636938 -4618 637174
rect -4534 636938 -4298 637174
rect -4854 636618 -4618 636854
rect -4534 636618 -4298 636854
rect -4854 600938 -4618 601174
rect -4534 600938 -4298 601174
rect -4854 600618 -4618 600854
rect -4534 600618 -4298 600854
rect -4854 564938 -4618 565174
rect -4534 564938 -4298 565174
rect -4854 564618 -4618 564854
rect -4534 564618 -4298 564854
rect -4854 528938 -4618 529174
rect -4534 528938 -4298 529174
rect -4854 528618 -4618 528854
rect -4534 528618 -4298 528854
rect -4854 492938 -4618 493174
rect -4534 492938 -4298 493174
rect -4854 492618 -4618 492854
rect -4534 492618 -4298 492854
rect -4854 456938 -4618 457174
rect -4534 456938 -4298 457174
rect -4854 456618 -4618 456854
rect -4534 456618 -4298 456854
rect -4854 420938 -4618 421174
rect -4534 420938 -4298 421174
rect -4854 420618 -4618 420854
rect -4534 420618 -4298 420854
rect -4854 384938 -4618 385174
rect -4534 384938 -4298 385174
rect -4854 384618 -4618 384854
rect -4534 384618 -4298 384854
rect -4854 348938 -4618 349174
rect -4534 348938 -4298 349174
rect -4854 348618 -4618 348854
rect -4534 348618 -4298 348854
rect -4854 312938 -4618 313174
rect -4534 312938 -4298 313174
rect -4854 312618 -4618 312854
rect -4534 312618 -4298 312854
rect -4854 276938 -4618 277174
rect -4534 276938 -4298 277174
rect -4854 276618 -4618 276854
rect -4534 276618 -4298 276854
rect -4854 240938 -4618 241174
rect -4534 240938 -4298 241174
rect -4854 240618 -4618 240854
rect -4534 240618 -4298 240854
rect -4854 204938 -4618 205174
rect -4534 204938 -4298 205174
rect -4854 204618 -4618 204854
rect -4534 204618 -4298 204854
rect -4854 168938 -4618 169174
rect -4534 168938 -4298 169174
rect -4854 168618 -4618 168854
rect -4534 168618 -4298 168854
rect -4854 132938 -4618 133174
rect -4534 132938 -4298 133174
rect -4854 132618 -4618 132854
rect -4534 132618 -4298 132854
rect -4854 96938 -4618 97174
rect -4534 96938 -4298 97174
rect -4854 96618 -4618 96854
rect -4534 96618 -4298 96854
rect -4854 60938 -4618 61174
rect -4534 60938 -4298 61174
rect -4854 60618 -4618 60854
rect -4534 60618 -4298 60854
rect -4854 24938 -4618 25174
rect -4534 24938 -4298 25174
rect -4854 24618 -4618 24854
rect -4534 24618 -4298 24854
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect 5546 706522 5782 706758
rect 5866 706522 6102 706758
rect 5546 706202 5782 706438
rect 5866 706202 6102 706438
rect -3894 690938 -3658 691174
rect -3574 690938 -3338 691174
rect -3894 690618 -3658 690854
rect -3574 690618 -3338 690854
rect -3894 654938 -3658 655174
rect -3574 654938 -3338 655174
rect -3894 654618 -3658 654854
rect -3574 654618 -3338 654854
rect -3894 618938 -3658 619174
rect -3574 618938 -3338 619174
rect -3894 618618 -3658 618854
rect -3574 618618 -3338 618854
rect -3894 582938 -3658 583174
rect -3574 582938 -3338 583174
rect -3894 582618 -3658 582854
rect -3574 582618 -3338 582854
rect -3894 546938 -3658 547174
rect -3574 546938 -3338 547174
rect -3894 546618 -3658 546854
rect -3574 546618 -3338 546854
rect -3894 510938 -3658 511174
rect -3574 510938 -3338 511174
rect -3894 510618 -3658 510854
rect -3574 510618 -3338 510854
rect -3894 474938 -3658 475174
rect -3574 474938 -3338 475174
rect -3894 474618 -3658 474854
rect -3574 474618 -3338 474854
rect -3894 438938 -3658 439174
rect -3574 438938 -3338 439174
rect -3894 438618 -3658 438854
rect -3574 438618 -3338 438854
rect -3894 402938 -3658 403174
rect -3574 402938 -3338 403174
rect -3894 402618 -3658 402854
rect -3574 402618 -3338 402854
rect -3894 366938 -3658 367174
rect -3574 366938 -3338 367174
rect -3894 366618 -3658 366854
rect -3574 366618 -3338 366854
rect -3894 330938 -3658 331174
rect -3574 330938 -3338 331174
rect -3894 330618 -3658 330854
rect -3574 330618 -3338 330854
rect -3894 294938 -3658 295174
rect -3574 294938 -3338 295174
rect -3894 294618 -3658 294854
rect -3574 294618 -3338 294854
rect -3894 258938 -3658 259174
rect -3574 258938 -3338 259174
rect -3894 258618 -3658 258854
rect -3574 258618 -3338 258854
rect -3894 222938 -3658 223174
rect -3574 222938 -3338 223174
rect -3894 222618 -3658 222854
rect -3574 222618 -3338 222854
rect -3894 186938 -3658 187174
rect -3574 186938 -3338 187174
rect -3894 186618 -3658 186854
rect -3574 186618 -3338 186854
rect -3894 150938 -3658 151174
rect -3574 150938 -3338 151174
rect -3894 150618 -3658 150854
rect -3574 150618 -3338 150854
rect -3894 114938 -3658 115174
rect -3574 114938 -3338 115174
rect -3894 114618 -3658 114854
rect -3574 114618 -3338 114854
rect -3894 78938 -3658 79174
rect -3574 78938 -3338 79174
rect -3894 78618 -3658 78854
rect -3574 78618 -3338 78854
rect -3894 42938 -3658 43174
rect -3574 42938 -3338 43174
rect -3894 42618 -3658 42854
rect -3574 42618 -3338 42854
rect -3894 6938 -3658 7174
rect -3574 6938 -3338 7174
rect -3894 6618 -3658 6854
rect -3574 6618 -3338 6854
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 669218 -2698 669454
rect -2614 669218 -2378 669454
rect -2934 668898 -2698 669134
rect -2614 668898 -2378 669134
rect -2934 633218 -2698 633454
rect -2614 633218 -2378 633454
rect -2934 632898 -2698 633134
rect -2614 632898 -2378 633134
rect -2934 597218 -2698 597454
rect -2614 597218 -2378 597454
rect -2934 596898 -2698 597134
rect -2614 596898 -2378 597134
rect -2934 561218 -2698 561454
rect -2614 561218 -2378 561454
rect -2934 560898 -2698 561134
rect -2614 560898 -2378 561134
rect -2934 525218 -2698 525454
rect -2614 525218 -2378 525454
rect -2934 524898 -2698 525134
rect -2614 524898 -2378 525134
rect -2934 489218 -2698 489454
rect -2614 489218 -2378 489454
rect -2934 488898 -2698 489134
rect -2614 488898 -2378 489134
rect -2934 453218 -2698 453454
rect -2614 453218 -2378 453454
rect -2934 452898 -2698 453134
rect -2614 452898 -2378 453134
rect -2934 417218 -2698 417454
rect -2614 417218 -2378 417454
rect -2934 416898 -2698 417134
rect -2614 416898 -2378 417134
rect -2934 381218 -2698 381454
rect -2614 381218 -2378 381454
rect -2934 380898 -2698 381134
rect -2614 380898 -2378 381134
rect -2934 345218 -2698 345454
rect -2614 345218 -2378 345454
rect -2934 344898 -2698 345134
rect -2614 344898 -2378 345134
rect -2934 309218 -2698 309454
rect -2614 309218 -2378 309454
rect -2934 308898 -2698 309134
rect -2614 308898 -2378 309134
rect -2934 273218 -2698 273454
rect -2614 273218 -2378 273454
rect -2934 272898 -2698 273134
rect -2614 272898 -2378 273134
rect -2934 237218 -2698 237454
rect -2614 237218 -2378 237454
rect -2934 236898 -2698 237134
rect -2614 236898 -2378 237134
rect -2934 201218 -2698 201454
rect -2614 201218 -2378 201454
rect -2934 200898 -2698 201134
rect -2614 200898 -2378 201134
rect -2934 165218 -2698 165454
rect -2614 165218 -2378 165454
rect -2934 164898 -2698 165134
rect -2614 164898 -2378 165134
rect -2934 129218 -2698 129454
rect -2614 129218 -2378 129454
rect -2934 128898 -2698 129134
rect -2614 128898 -2378 129134
rect -2934 93218 -2698 93454
rect -2614 93218 -2378 93454
rect -2934 92898 -2698 93134
rect -2614 92898 -2378 93134
rect -2934 57218 -2698 57454
rect -2614 57218 -2378 57454
rect -2934 56898 -2698 57134
rect -2614 56898 -2378 57134
rect -2934 21218 -2698 21454
rect -2614 21218 -2378 21454
rect -2934 20898 -2698 21134
rect -2614 20898 -2378 21134
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect 5546 -2502 5782 -2266
rect 5866 -2502 6102 -2266
rect 5546 -2822 5782 -2586
rect 5866 -2822 6102 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 9266 658658 9502 658894
rect 9586 658658 9822 658894
rect 9266 658338 9502 658574
rect 9586 658338 9822 658574
rect 9266 622658 9502 622894
rect 9586 622658 9822 622894
rect 9266 622338 9502 622574
rect 9586 622338 9822 622574
rect 9266 586658 9502 586894
rect 9586 586658 9822 586894
rect 9266 586338 9502 586574
rect 9586 586338 9822 586574
rect 9266 550658 9502 550894
rect 9586 550658 9822 550894
rect 9266 550338 9502 550574
rect 9586 550338 9822 550574
rect 9266 514658 9502 514894
rect 9586 514658 9822 514894
rect 9266 514338 9502 514574
rect 9586 514338 9822 514574
rect 9266 478658 9502 478894
rect 9586 478658 9822 478894
rect 9266 478338 9502 478574
rect 9586 478338 9822 478574
rect 9266 442658 9502 442894
rect 9586 442658 9822 442894
rect 9266 442338 9502 442574
rect 9586 442338 9822 442574
rect 9266 406658 9502 406894
rect 9586 406658 9822 406894
rect 9266 406338 9502 406574
rect 9586 406338 9822 406574
rect 9266 370658 9502 370894
rect 9586 370658 9822 370894
rect 9266 370338 9502 370574
rect 9586 370338 9822 370574
rect 9266 334658 9502 334894
rect 9586 334658 9822 334894
rect 9266 334338 9502 334574
rect 9586 334338 9822 334574
rect 9266 298658 9502 298894
rect 9586 298658 9822 298894
rect 9266 298338 9502 298574
rect 9586 298338 9822 298574
rect 9266 262658 9502 262894
rect 9586 262658 9822 262894
rect 9266 262338 9502 262574
rect 9586 262338 9822 262574
rect 9266 226658 9502 226894
rect 9586 226658 9822 226894
rect 9266 226338 9502 226574
rect 9586 226338 9822 226574
rect 9266 190658 9502 190894
rect 9586 190658 9822 190894
rect 9266 190338 9502 190574
rect 9586 190338 9822 190574
rect 9266 154658 9502 154894
rect 9586 154658 9822 154894
rect 9266 154338 9502 154574
rect 9586 154338 9822 154574
rect 9266 118658 9502 118894
rect 9586 118658 9822 118894
rect 9266 118338 9502 118574
rect 9586 118338 9822 118574
rect 9266 82658 9502 82894
rect 9586 82658 9822 82894
rect 9266 82338 9502 82574
rect 9586 82338 9822 82574
rect 9266 46658 9502 46894
rect 9586 46658 9822 46894
rect 9266 46338 9502 46574
rect 9586 46338 9822 46574
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect 9266 -4422 9502 -4186
rect 9586 -4422 9822 -4186
rect 9266 -4742 9502 -4506
rect 9586 -4742 9822 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect 30986 711322 31222 711558
rect 31306 711322 31542 711558
rect 30986 711002 31222 711238
rect 31306 711002 31542 711238
rect 27266 709402 27502 709638
rect 27586 709402 27822 709638
rect 27266 709082 27502 709318
rect 27586 709082 27822 709318
rect 23546 707482 23782 707718
rect 23866 707482 24102 707718
rect 23546 707162 23782 707398
rect 23866 707162 24102 707398
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 12986 662378 13222 662614
rect 13306 662378 13542 662614
rect 12986 662058 13222 662294
rect 13306 662058 13542 662294
rect 12986 626378 13222 626614
rect 13306 626378 13542 626614
rect 12986 626058 13222 626294
rect 13306 626058 13542 626294
rect 12986 590378 13222 590614
rect 13306 590378 13542 590614
rect 12986 590058 13222 590294
rect 13306 590058 13542 590294
rect 12986 554378 13222 554614
rect 13306 554378 13542 554614
rect 12986 554058 13222 554294
rect 13306 554058 13542 554294
rect 12986 518378 13222 518614
rect 13306 518378 13542 518614
rect 12986 518058 13222 518294
rect 13306 518058 13542 518294
rect 12986 482378 13222 482614
rect 13306 482378 13542 482614
rect 12986 482058 13222 482294
rect 13306 482058 13542 482294
rect 12986 446378 13222 446614
rect 13306 446378 13542 446614
rect 12986 446058 13222 446294
rect 13306 446058 13542 446294
rect 12986 410378 13222 410614
rect 13306 410378 13542 410614
rect 12986 410058 13222 410294
rect 13306 410058 13542 410294
rect 12986 374378 13222 374614
rect 13306 374378 13542 374614
rect 12986 374058 13222 374294
rect 13306 374058 13542 374294
rect 12986 338378 13222 338614
rect 13306 338378 13542 338614
rect 12986 338058 13222 338294
rect 13306 338058 13542 338294
rect 12986 302378 13222 302614
rect 13306 302378 13542 302614
rect 12986 302058 13222 302294
rect 13306 302058 13542 302294
rect 12986 266378 13222 266614
rect 13306 266378 13542 266614
rect 12986 266058 13222 266294
rect 13306 266058 13542 266294
rect 12986 230378 13222 230614
rect 13306 230378 13542 230614
rect 12986 230058 13222 230294
rect 13306 230058 13542 230294
rect 12986 194378 13222 194614
rect 13306 194378 13542 194614
rect 12986 194058 13222 194294
rect 13306 194058 13542 194294
rect 12986 158378 13222 158614
rect 13306 158378 13542 158614
rect 12986 158058 13222 158294
rect 13306 158058 13542 158294
rect 12986 122378 13222 122614
rect 13306 122378 13542 122614
rect 12986 122058 13222 122294
rect 13306 122058 13542 122294
rect 12986 86378 13222 86614
rect 13306 86378 13542 86614
rect 12986 86058 13222 86294
rect 13306 86058 13542 86294
rect 12986 50378 13222 50614
rect 13306 50378 13542 50614
rect 12986 50058 13222 50294
rect 13306 50058 13542 50294
rect 12986 14378 13222 14614
rect 13306 14378 13542 14614
rect 12986 14058 13222 14294
rect 13306 14058 13542 14294
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect 19826 705562 20062 705798
rect 20146 705562 20382 705798
rect 19826 705242 20062 705478
rect 20146 705242 20382 705478
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -1542 20062 -1306
rect 20146 -1542 20382 -1306
rect 19826 -1862 20062 -1626
rect 20146 -1862 20382 -1626
rect 23546 672938 23782 673174
rect 23866 672938 24102 673174
rect 23546 672618 23782 672854
rect 23866 672618 24102 672854
rect 23546 636938 23782 637174
rect 23866 636938 24102 637174
rect 23546 636618 23782 636854
rect 23866 636618 24102 636854
rect 23546 600938 23782 601174
rect 23866 600938 24102 601174
rect 23546 600618 23782 600854
rect 23866 600618 24102 600854
rect 23546 564938 23782 565174
rect 23866 564938 24102 565174
rect 23546 564618 23782 564854
rect 23866 564618 24102 564854
rect 23546 528938 23782 529174
rect 23866 528938 24102 529174
rect 23546 528618 23782 528854
rect 23866 528618 24102 528854
rect 23546 492938 23782 493174
rect 23866 492938 24102 493174
rect 23546 492618 23782 492854
rect 23866 492618 24102 492854
rect 23546 456938 23782 457174
rect 23866 456938 24102 457174
rect 23546 456618 23782 456854
rect 23866 456618 24102 456854
rect 23546 420938 23782 421174
rect 23866 420938 24102 421174
rect 23546 420618 23782 420854
rect 23866 420618 24102 420854
rect 23546 384938 23782 385174
rect 23866 384938 24102 385174
rect 23546 384618 23782 384854
rect 23866 384618 24102 384854
rect 23546 348938 23782 349174
rect 23866 348938 24102 349174
rect 23546 348618 23782 348854
rect 23866 348618 24102 348854
rect 23546 312938 23782 313174
rect 23866 312938 24102 313174
rect 23546 312618 23782 312854
rect 23866 312618 24102 312854
rect 23546 276938 23782 277174
rect 23866 276938 24102 277174
rect 23546 276618 23782 276854
rect 23866 276618 24102 276854
rect 23546 240938 23782 241174
rect 23866 240938 24102 241174
rect 23546 240618 23782 240854
rect 23866 240618 24102 240854
rect 23546 204938 23782 205174
rect 23866 204938 24102 205174
rect 23546 204618 23782 204854
rect 23866 204618 24102 204854
rect 23546 168938 23782 169174
rect 23866 168938 24102 169174
rect 23546 168618 23782 168854
rect 23866 168618 24102 168854
rect 23546 132938 23782 133174
rect 23866 132938 24102 133174
rect 23546 132618 23782 132854
rect 23866 132618 24102 132854
rect 23546 96938 23782 97174
rect 23866 96938 24102 97174
rect 23546 96618 23782 96854
rect 23866 96618 24102 96854
rect 23546 60938 23782 61174
rect 23866 60938 24102 61174
rect 23546 60618 23782 60854
rect 23866 60618 24102 60854
rect 23546 24938 23782 25174
rect 23866 24938 24102 25174
rect 23546 24618 23782 24854
rect 23866 24618 24102 24854
rect 23546 -3462 23782 -3226
rect 23866 -3462 24102 -3226
rect 23546 -3782 23782 -3546
rect 23866 -3782 24102 -3546
rect 27266 676658 27502 676894
rect 27586 676658 27822 676894
rect 27266 676338 27502 676574
rect 27586 676338 27822 676574
rect 27266 640658 27502 640894
rect 27586 640658 27822 640894
rect 27266 640338 27502 640574
rect 27586 640338 27822 640574
rect 27266 604658 27502 604894
rect 27586 604658 27822 604894
rect 27266 604338 27502 604574
rect 27586 604338 27822 604574
rect 27266 568658 27502 568894
rect 27586 568658 27822 568894
rect 27266 568338 27502 568574
rect 27586 568338 27822 568574
rect 27266 532658 27502 532894
rect 27586 532658 27822 532894
rect 27266 532338 27502 532574
rect 27586 532338 27822 532574
rect 27266 496658 27502 496894
rect 27586 496658 27822 496894
rect 27266 496338 27502 496574
rect 27586 496338 27822 496574
rect 27266 460658 27502 460894
rect 27586 460658 27822 460894
rect 27266 460338 27502 460574
rect 27586 460338 27822 460574
rect 27266 424658 27502 424894
rect 27586 424658 27822 424894
rect 27266 424338 27502 424574
rect 27586 424338 27822 424574
rect 27266 388658 27502 388894
rect 27586 388658 27822 388894
rect 27266 388338 27502 388574
rect 27586 388338 27822 388574
rect 27266 352658 27502 352894
rect 27586 352658 27822 352894
rect 27266 352338 27502 352574
rect 27586 352338 27822 352574
rect 27266 316658 27502 316894
rect 27586 316658 27822 316894
rect 27266 316338 27502 316574
rect 27586 316338 27822 316574
rect 27266 280658 27502 280894
rect 27586 280658 27822 280894
rect 27266 280338 27502 280574
rect 27586 280338 27822 280574
rect 27266 244658 27502 244894
rect 27586 244658 27822 244894
rect 27266 244338 27502 244574
rect 27586 244338 27822 244574
rect 27266 208658 27502 208894
rect 27586 208658 27822 208894
rect 27266 208338 27502 208574
rect 27586 208338 27822 208574
rect 27266 172658 27502 172894
rect 27586 172658 27822 172894
rect 27266 172338 27502 172574
rect 27586 172338 27822 172574
rect 27266 136658 27502 136894
rect 27586 136658 27822 136894
rect 27266 136338 27502 136574
rect 27586 136338 27822 136574
rect 27266 100658 27502 100894
rect 27586 100658 27822 100894
rect 27266 100338 27502 100574
rect 27586 100338 27822 100574
rect 27266 64658 27502 64894
rect 27586 64658 27822 64894
rect 27266 64338 27502 64574
rect 27586 64338 27822 64574
rect 27266 28658 27502 28894
rect 27586 28658 27822 28894
rect 27266 28338 27502 28574
rect 27586 28338 27822 28574
rect 27266 -5382 27502 -5146
rect 27586 -5382 27822 -5146
rect 27266 -5702 27502 -5466
rect 27586 -5702 27822 -5466
rect 48986 710362 49222 710598
rect 49306 710362 49542 710598
rect 48986 710042 49222 710278
rect 49306 710042 49542 710278
rect 45266 708442 45502 708678
rect 45586 708442 45822 708678
rect 45266 708122 45502 708358
rect 45586 708122 45822 708358
rect 41546 706522 41782 706758
rect 41866 706522 42102 706758
rect 41546 706202 41782 706438
rect 41866 706202 42102 706438
rect 30986 680378 31222 680614
rect 31306 680378 31542 680614
rect 30986 680058 31222 680294
rect 31306 680058 31542 680294
rect 30986 644378 31222 644614
rect 31306 644378 31542 644614
rect 30986 644058 31222 644294
rect 31306 644058 31542 644294
rect 30986 608378 31222 608614
rect 31306 608378 31542 608614
rect 30986 608058 31222 608294
rect 31306 608058 31542 608294
rect 30986 572378 31222 572614
rect 31306 572378 31542 572614
rect 30986 572058 31222 572294
rect 31306 572058 31542 572294
rect 30986 536378 31222 536614
rect 31306 536378 31542 536614
rect 30986 536058 31222 536294
rect 31306 536058 31542 536294
rect 30986 500378 31222 500614
rect 31306 500378 31542 500614
rect 30986 500058 31222 500294
rect 31306 500058 31542 500294
rect 30986 464378 31222 464614
rect 31306 464378 31542 464614
rect 30986 464058 31222 464294
rect 31306 464058 31542 464294
rect 30986 428378 31222 428614
rect 31306 428378 31542 428614
rect 30986 428058 31222 428294
rect 31306 428058 31542 428294
rect 30986 392378 31222 392614
rect 31306 392378 31542 392614
rect 30986 392058 31222 392294
rect 31306 392058 31542 392294
rect 30986 356378 31222 356614
rect 31306 356378 31542 356614
rect 30986 356058 31222 356294
rect 31306 356058 31542 356294
rect 30986 320378 31222 320614
rect 31306 320378 31542 320614
rect 30986 320058 31222 320294
rect 31306 320058 31542 320294
rect 30986 284378 31222 284614
rect 31306 284378 31542 284614
rect 30986 284058 31222 284294
rect 31306 284058 31542 284294
rect 30986 248378 31222 248614
rect 31306 248378 31542 248614
rect 30986 248058 31222 248294
rect 31306 248058 31542 248294
rect 30986 212378 31222 212614
rect 31306 212378 31542 212614
rect 30986 212058 31222 212294
rect 31306 212058 31542 212294
rect 30986 176378 31222 176614
rect 31306 176378 31542 176614
rect 30986 176058 31222 176294
rect 31306 176058 31542 176294
rect 30986 140378 31222 140614
rect 31306 140378 31542 140614
rect 30986 140058 31222 140294
rect 31306 140058 31542 140294
rect 30986 104378 31222 104614
rect 31306 104378 31542 104614
rect 30986 104058 31222 104294
rect 31306 104058 31542 104294
rect 30986 68378 31222 68614
rect 31306 68378 31542 68614
rect 30986 68058 31222 68294
rect 31306 68058 31542 68294
rect 30986 32378 31222 32614
rect 31306 32378 31542 32614
rect 30986 32058 31222 32294
rect 31306 32058 31542 32294
rect 12986 -6342 13222 -6106
rect 13306 -6342 13542 -6106
rect 12986 -6662 13222 -6426
rect 13306 -6662 13542 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 41546 654938 41782 655174
rect 41866 654938 42102 655174
rect 41546 654618 41782 654854
rect 41866 654618 42102 654854
rect 41546 618938 41782 619174
rect 41866 618938 42102 619174
rect 41546 618618 41782 618854
rect 41866 618618 42102 618854
rect 41546 582938 41782 583174
rect 41866 582938 42102 583174
rect 41546 582618 41782 582854
rect 41866 582618 42102 582854
rect 41546 546938 41782 547174
rect 41866 546938 42102 547174
rect 41546 546618 41782 546854
rect 41866 546618 42102 546854
rect 41546 510938 41782 511174
rect 41866 510938 42102 511174
rect 41546 510618 41782 510854
rect 41866 510618 42102 510854
rect 41546 474938 41782 475174
rect 41866 474938 42102 475174
rect 41546 474618 41782 474854
rect 41866 474618 42102 474854
rect 41546 438938 41782 439174
rect 41866 438938 42102 439174
rect 41546 438618 41782 438854
rect 41866 438618 42102 438854
rect 41546 402938 41782 403174
rect 41866 402938 42102 403174
rect 41546 402618 41782 402854
rect 41866 402618 42102 402854
rect 41546 366938 41782 367174
rect 41866 366938 42102 367174
rect 41546 366618 41782 366854
rect 41866 366618 42102 366854
rect 41546 330938 41782 331174
rect 41866 330938 42102 331174
rect 41546 330618 41782 330854
rect 41866 330618 42102 330854
rect 41546 294938 41782 295174
rect 41866 294938 42102 295174
rect 41546 294618 41782 294854
rect 41866 294618 42102 294854
rect 41546 258938 41782 259174
rect 41866 258938 42102 259174
rect 41546 258618 41782 258854
rect 41866 258618 42102 258854
rect 41546 222938 41782 223174
rect 41866 222938 42102 223174
rect 41546 222618 41782 222854
rect 41866 222618 42102 222854
rect 41546 186938 41782 187174
rect 41866 186938 42102 187174
rect 41546 186618 41782 186854
rect 41866 186618 42102 186854
rect 41546 150938 41782 151174
rect 41866 150938 42102 151174
rect 41546 150618 41782 150854
rect 41866 150618 42102 150854
rect 41546 114938 41782 115174
rect 41866 114938 42102 115174
rect 41546 114618 41782 114854
rect 41866 114618 42102 114854
rect 41546 78938 41782 79174
rect 41866 78938 42102 79174
rect 41546 78618 41782 78854
rect 41866 78618 42102 78854
rect 41546 42938 41782 43174
rect 41866 42938 42102 43174
rect 41546 42618 41782 42854
rect 41866 42618 42102 42854
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -2502 41782 -2266
rect 41866 -2502 42102 -2266
rect 41546 -2822 41782 -2586
rect 41866 -2822 42102 -2586
rect 45266 694658 45502 694894
rect 45586 694658 45822 694894
rect 45266 694338 45502 694574
rect 45586 694338 45822 694574
rect 45266 658658 45502 658894
rect 45586 658658 45822 658894
rect 45266 658338 45502 658574
rect 45586 658338 45822 658574
rect 45266 622658 45502 622894
rect 45586 622658 45822 622894
rect 45266 622338 45502 622574
rect 45586 622338 45822 622574
rect 45266 586658 45502 586894
rect 45586 586658 45822 586894
rect 45266 586338 45502 586574
rect 45586 586338 45822 586574
rect 45266 550658 45502 550894
rect 45586 550658 45822 550894
rect 45266 550338 45502 550574
rect 45586 550338 45822 550574
rect 45266 514658 45502 514894
rect 45586 514658 45822 514894
rect 45266 514338 45502 514574
rect 45586 514338 45822 514574
rect 45266 478658 45502 478894
rect 45586 478658 45822 478894
rect 45266 478338 45502 478574
rect 45586 478338 45822 478574
rect 66986 711322 67222 711558
rect 67306 711322 67542 711558
rect 66986 711002 67222 711238
rect 67306 711002 67542 711238
rect 63266 709402 63502 709638
rect 63586 709402 63822 709638
rect 63266 709082 63502 709318
rect 63586 709082 63822 709318
rect 59546 707482 59782 707718
rect 59866 707482 60102 707718
rect 59546 707162 59782 707398
rect 59866 707162 60102 707398
rect 48986 698378 49222 698614
rect 49306 698378 49542 698614
rect 48986 698058 49222 698294
rect 49306 698058 49542 698294
rect 48986 662378 49222 662614
rect 49306 662378 49542 662614
rect 48986 662058 49222 662294
rect 49306 662058 49542 662294
rect 48986 626378 49222 626614
rect 49306 626378 49542 626614
rect 48986 626058 49222 626294
rect 49306 626058 49542 626294
rect 48986 590378 49222 590614
rect 49306 590378 49542 590614
rect 48986 590058 49222 590294
rect 49306 590058 49542 590294
rect 48986 554378 49222 554614
rect 49306 554378 49542 554614
rect 48986 554058 49222 554294
rect 49306 554058 49542 554294
rect 48986 518378 49222 518614
rect 49306 518378 49542 518614
rect 48986 518058 49222 518294
rect 49306 518058 49542 518294
rect 48986 482378 49222 482614
rect 49306 482378 49542 482614
rect 48986 482058 49222 482294
rect 49306 482058 49542 482294
rect 55826 705562 56062 705798
rect 56146 705562 56382 705798
rect 55826 705242 56062 705478
rect 56146 705242 56382 705478
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 59546 672938 59782 673174
rect 59866 672938 60102 673174
rect 59546 672618 59782 672854
rect 59866 672618 60102 672854
rect 59546 636938 59782 637174
rect 59866 636938 60102 637174
rect 59546 636618 59782 636854
rect 59866 636618 60102 636854
rect 59546 600938 59782 601174
rect 59866 600938 60102 601174
rect 59546 600618 59782 600854
rect 59866 600618 60102 600854
rect 59546 564938 59782 565174
rect 59866 564938 60102 565174
rect 59546 564618 59782 564854
rect 59866 564618 60102 564854
rect 59546 528938 59782 529174
rect 59866 528938 60102 529174
rect 59546 528618 59782 528854
rect 59866 528618 60102 528854
rect 59546 492938 59782 493174
rect 59866 492938 60102 493174
rect 59546 492618 59782 492854
rect 59866 492618 60102 492854
rect 63266 676658 63502 676894
rect 63586 676658 63822 676894
rect 63266 676338 63502 676574
rect 63586 676338 63822 676574
rect 63266 640658 63502 640894
rect 63586 640658 63822 640894
rect 63266 640338 63502 640574
rect 63586 640338 63822 640574
rect 63266 604658 63502 604894
rect 63586 604658 63822 604894
rect 63266 604338 63502 604574
rect 63586 604338 63822 604574
rect 63266 568658 63502 568894
rect 63586 568658 63822 568894
rect 63266 568338 63502 568574
rect 63586 568338 63822 568574
rect 63266 532658 63502 532894
rect 63586 532658 63822 532894
rect 63266 532338 63502 532574
rect 63586 532338 63822 532574
rect 63266 496658 63502 496894
rect 63586 496658 63822 496894
rect 63266 496338 63502 496574
rect 63586 496338 63822 496574
rect 84986 710362 85222 710598
rect 85306 710362 85542 710598
rect 84986 710042 85222 710278
rect 85306 710042 85542 710278
rect 81266 708442 81502 708678
rect 81586 708442 81822 708678
rect 81266 708122 81502 708358
rect 81586 708122 81822 708358
rect 77546 706522 77782 706758
rect 77866 706522 78102 706758
rect 77546 706202 77782 706438
rect 77866 706202 78102 706438
rect 66986 680378 67222 680614
rect 67306 680378 67542 680614
rect 66986 680058 67222 680294
rect 67306 680058 67542 680294
rect 66986 644378 67222 644614
rect 67306 644378 67542 644614
rect 66986 644058 67222 644294
rect 67306 644058 67542 644294
rect 66986 608378 67222 608614
rect 67306 608378 67542 608614
rect 66986 608058 67222 608294
rect 67306 608058 67542 608294
rect 66986 572378 67222 572614
rect 67306 572378 67542 572614
rect 66986 572058 67222 572294
rect 67306 572058 67542 572294
rect 66986 536378 67222 536614
rect 67306 536378 67542 536614
rect 66986 536058 67222 536294
rect 67306 536058 67542 536294
rect 66986 500378 67222 500614
rect 67306 500378 67542 500614
rect 66986 500058 67222 500294
rect 67306 500058 67542 500294
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 73826 579218 74062 579454
rect 74146 579218 74382 579454
rect 73826 578898 74062 579134
rect 74146 578898 74382 579134
rect 73826 543218 74062 543454
rect 74146 543218 74382 543454
rect 73826 542898 74062 543134
rect 74146 542898 74382 543134
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 77546 654938 77782 655174
rect 77866 654938 78102 655174
rect 77546 654618 77782 654854
rect 77866 654618 78102 654854
rect 77546 618938 77782 619174
rect 77866 618938 78102 619174
rect 77546 618618 77782 618854
rect 77866 618618 78102 618854
rect 77546 582938 77782 583174
rect 77866 582938 78102 583174
rect 77546 582618 77782 582854
rect 77866 582618 78102 582854
rect 77546 546938 77782 547174
rect 77866 546938 78102 547174
rect 77546 546618 77782 546854
rect 77866 546618 78102 546854
rect 77546 510938 77782 511174
rect 77866 510938 78102 511174
rect 77546 510618 77782 510854
rect 77866 510618 78102 510854
rect 77546 474938 77782 475174
rect 77866 474938 78102 475174
rect 77546 474618 77782 474854
rect 77866 474618 78102 474854
rect 81266 694658 81502 694894
rect 81586 694658 81822 694894
rect 81266 694338 81502 694574
rect 81586 694338 81822 694574
rect 81266 658658 81502 658894
rect 81586 658658 81822 658894
rect 81266 658338 81502 658574
rect 81586 658338 81822 658574
rect 81266 622658 81502 622894
rect 81586 622658 81822 622894
rect 81266 622338 81502 622574
rect 81586 622338 81822 622574
rect 81266 586658 81502 586894
rect 81586 586658 81822 586894
rect 81266 586338 81502 586574
rect 81586 586338 81822 586574
rect 81266 550658 81502 550894
rect 81586 550658 81822 550894
rect 81266 550338 81502 550574
rect 81586 550338 81822 550574
rect 81266 514658 81502 514894
rect 81586 514658 81822 514894
rect 81266 514338 81502 514574
rect 81586 514338 81822 514574
rect 81266 478658 81502 478894
rect 81586 478658 81822 478894
rect 81266 478338 81502 478574
rect 81586 478338 81822 478574
rect 102986 711322 103222 711558
rect 103306 711322 103542 711558
rect 102986 711002 103222 711238
rect 103306 711002 103542 711238
rect 99266 709402 99502 709638
rect 99586 709402 99822 709638
rect 99266 709082 99502 709318
rect 99586 709082 99822 709318
rect 95546 707482 95782 707718
rect 95866 707482 96102 707718
rect 95546 707162 95782 707398
rect 95866 707162 96102 707398
rect 84986 698378 85222 698614
rect 85306 698378 85542 698614
rect 84986 698058 85222 698294
rect 85306 698058 85542 698294
rect 84986 662378 85222 662614
rect 85306 662378 85542 662614
rect 84986 662058 85222 662294
rect 85306 662058 85542 662294
rect 84986 626378 85222 626614
rect 85306 626378 85542 626614
rect 84986 626058 85222 626294
rect 85306 626058 85542 626294
rect 84986 590378 85222 590614
rect 85306 590378 85542 590614
rect 84986 590058 85222 590294
rect 85306 590058 85542 590294
rect 84986 554378 85222 554614
rect 85306 554378 85542 554614
rect 84986 554058 85222 554294
rect 85306 554058 85542 554294
rect 84986 518378 85222 518614
rect 85306 518378 85542 518614
rect 84986 518058 85222 518294
rect 85306 518058 85542 518294
rect 84986 482378 85222 482614
rect 85306 482378 85542 482614
rect 84986 482058 85222 482294
rect 85306 482058 85542 482294
rect 91826 705562 92062 705798
rect 92146 705562 92382 705798
rect 91826 705242 92062 705478
rect 92146 705242 92382 705478
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 91826 561218 92062 561454
rect 92146 561218 92382 561454
rect 91826 560898 92062 561134
rect 92146 560898 92382 561134
rect 91826 525218 92062 525454
rect 92146 525218 92382 525454
rect 91826 524898 92062 525134
rect 92146 524898 92382 525134
rect 91826 489218 92062 489454
rect 92146 489218 92382 489454
rect 91826 488898 92062 489134
rect 92146 488898 92382 489134
rect 95546 672938 95782 673174
rect 95866 672938 96102 673174
rect 95546 672618 95782 672854
rect 95866 672618 96102 672854
rect 95546 636938 95782 637174
rect 95866 636938 96102 637174
rect 95546 636618 95782 636854
rect 95866 636618 96102 636854
rect 95546 600938 95782 601174
rect 95866 600938 96102 601174
rect 95546 600618 95782 600854
rect 95866 600618 96102 600854
rect 95546 564938 95782 565174
rect 95866 564938 96102 565174
rect 95546 564618 95782 564854
rect 95866 564618 96102 564854
rect 95546 528938 95782 529174
rect 95866 528938 96102 529174
rect 95546 528618 95782 528854
rect 95866 528618 96102 528854
rect 95546 492938 95782 493174
rect 95866 492938 96102 493174
rect 95546 492618 95782 492854
rect 95866 492618 96102 492854
rect 99266 676658 99502 676894
rect 99586 676658 99822 676894
rect 99266 676338 99502 676574
rect 99586 676338 99822 676574
rect 99266 640658 99502 640894
rect 99586 640658 99822 640894
rect 99266 640338 99502 640574
rect 99586 640338 99822 640574
rect 99266 604658 99502 604894
rect 99586 604658 99822 604894
rect 99266 604338 99502 604574
rect 99586 604338 99822 604574
rect 99266 568658 99502 568894
rect 99586 568658 99822 568894
rect 99266 568338 99502 568574
rect 99586 568338 99822 568574
rect 99266 532658 99502 532894
rect 99586 532658 99822 532894
rect 99266 532338 99502 532574
rect 99586 532338 99822 532574
rect 99266 496658 99502 496894
rect 99586 496658 99822 496894
rect 99266 496338 99502 496574
rect 99586 496338 99822 496574
rect 120986 710362 121222 710598
rect 121306 710362 121542 710598
rect 120986 710042 121222 710278
rect 121306 710042 121542 710278
rect 117266 708442 117502 708678
rect 117586 708442 117822 708678
rect 117266 708122 117502 708358
rect 117586 708122 117822 708358
rect 113546 706522 113782 706758
rect 113866 706522 114102 706758
rect 113546 706202 113782 706438
rect 113866 706202 114102 706438
rect 102986 680378 103222 680614
rect 103306 680378 103542 680614
rect 102986 680058 103222 680294
rect 103306 680058 103542 680294
rect 102986 644378 103222 644614
rect 103306 644378 103542 644614
rect 102986 644058 103222 644294
rect 103306 644058 103542 644294
rect 102986 608378 103222 608614
rect 103306 608378 103542 608614
rect 102986 608058 103222 608294
rect 103306 608058 103542 608294
rect 102986 572378 103222 572614
rect 103306 572378 103542 572614
rect 102986 572058 103222 572294
rect 103306 572058 103542 572294
rect 102986 536378 103222 536614
rect 103306 536378 103542 536614
rect 102986 536058 103222 536294
rect 103306 536058 103542 536294
rect 102986 500378 103222 500614
rect 103306 500378 103542 500614
rect 102986 500058 103222 500294
rect 103306 500058 103542 500294
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 109826 507218 110062 507454
rect 110146 507218 110382 507454
rect 109826 506898 110062 507134
rect 110146 506898 110382 507134
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 113546 654938 113782 655174
rect 113866 654938 114102 655174
rect 113546 654618 113782 654854
rect 113866 654618 114102 654854
rect 113546 618938 113782 619174
rect 113866 618938 114102 619174
rect 113546 618618 113782 618854
rect 113866 618618 114102 618854
rect 113546 582938 113782 583174
rect 113866 582938 114102 583174
rect 113546 582618 113782 582854
rect 113866 582618 114102 582854
rect 113546 546938 113782 547174
rect 113866 546938 114102 547174
rect 113546 546618 113782 546854
rect 113866 546618 114102 546854
rect 113546 510938 113782 511174
rect 113866 510938 114102 511174
rect 113546 510618 113782 510854
rect 113866 510618 114102 510854
rect 113546 474938 113782 475174
rect 113866 474938 114102 475174
rect 113546 474618 113782 474854
rect 113866 474618 114102 474854
rect 117266 694658 117502 694894
rect 117586 694658 117822 694894
rect 117266 694338 117502 694574
rect 117586 694338 117822 694574
rect 117266 658658 117502 658894
rect 117586 658658 117822 658894
rect 117266 658338 117502 658574
rect 117586 658338 117822 658574
rect 117266 622658 117502 622894
rect 117586 622658 117822 622894
rect 117266 622338 117502 622574
rect 117586 622338 117822 622574
rect 117266 586658 117502 586894
rect 117586 586658 117822 586894
rect 117266 586338 117502 586574
rect 117586 586338 117822 586574
rect 117266 550658 117502 550894
rect 117586 550658 117822 550894
rect 117266 550338 117502 550574
rect 117586 550338 117822 550574
rect 117266 514658 117502 514894
rect 117586 514658 117822 514894
rect 117266 514338 117502 514574
rect 117586 514338 117822 514574
rect 117266 478658 117502 478894
rect 117586 478658 117822 478894
rect 117266 478338 117502 478574
rect 117586 478338 117822 478574
rect 138986 711322 139222 711558
rect 139306 711322 139542 711558
rect 138986 711002 139222 711238
rect 139306 711002 139542 711238
rect 135266 709402 135502 709638
rect 135586 709402 135822 709638
rect 135266 709082 135502 709318
rect 135586 709082 135822 709318
rect 131546 707482 131782 707718
rect 131866 707482 132102 707718
rect 131546 707162 131782 707398
rect 131866 707162 132102 707398
rect 120986 698378 121222 698614
rect 121306 698378 121542 698614
rect 120986 698058 121222 698294
rect 121306 698058 121542 698294
rect 120986 662378 121222 662614
rect 121306 662378 121542 662614
rect 120986 662058 121222 662294
rect 121306 662058 121542 662294
rect 120986 626378 121222 626614
rect 121306 626378 121542 626614
rect 120986 626058 121222 626294
rect 121306 626058 121542 626294
rect 120986 590378 121222 590614
rect 121306 590378 121542 590614
rect 120986 590058 121222 590294
rect 121306 590058 121542 590294
rect 120986 554378 121222 554614
rect 121306 554378 121542 554614
rect 120986 554058 121222 554294
rect 121306 554058 121542 554294
rect 120986 518378 121222 518614
rect 121306 518378 121542 518614
rect 120986 518058 121222 518294
rect 121306 518058 121542 518294
rect 120986 482378 121222 482614
rect 121306 482378 121542 482614
rect 120986 482058 121222 482294
rect 121306 482058 121542 482294
rect 127826 705562 128062 705798
rect 128146 705562 128382 705798
rect 127826 705242 128062 705478
rect 128146 705242 128382 705478
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 127826 525218 128062 525454
rect 128146 525218 128382 525454
rect 127826 524898 128062 525134
rect 128146 524898 128382 525134
rect 127826 489218 128062 489454
rect 128146 489218 128382 489454
rect 127826 488898 128062 489134
rect 128146 488898 128382 489134
rect 131546 672938 131782 673174
rect 131866 672938 132102 673174
rect 131546 672618 131782 672854
rect 131866 672618 132102 672854
rect 131546 636938 131782 637174
rect 131866 636938 132102 637174
rect 131546 636618 131782 636854
rect 131866 636618 132102 636854
rect 131546 600938 131782 601174
rect 131866 600938 132102 601174
rect 131546 600618 131782 600854
rect 131866 600618 132102 600854
rect 131546 564938 131782 565174
rect 131866 564938 132102 565174
rect 131546 564618 131782 564854
rect 131866 564618 132102 564854
rect 131546 528938 131782 529174
rect 131866 528938 132102 529174
rect 131546 528618 131782 528854
rect 131866 528618 132102 528854
rect 131546 492938 131782 493174
rect 131866 492938 132102 493174
rect 131546 492618 131782 492854
rect 131866 492618 132102 492854
rect 135266 676658 135502 676894
rect 135586 676658 135822 676894
rect 135266 676338 135502 676574
rect 135586 676338 135822 676574
rect 135266 640658 135502 640894
rect 135586 640658 135822 640894
rect 135266 640338 135502 640574
rect 135586 640338 135822 640574
rect 135266 604658 135502 604894
rect 135586 604658 135822 604894
rect 135266 604338 135502 604574
rect 135586 604338 135822 604574
rect 135266 568658 135502 568894
rect 135586 568658 135822 568894
rect 135266 568338 135502 568574
rect 135586 568338 135822 568574
rect 135266 532658 135502 532894
rect 135586 532658 135822 532894
rect 135266 532338 135502 532574
rect 135586 532338 135822 532574
rect 135266 496658 135502 496894
rect 135586 496658 135822 496894
rect 135266 496338 135502 496574
rect 135586 496338 135822 496574
rect 156986 710362 157222 710598
rect 157306 710362 157542 710598
rect 156986 710042 157222 710278
rect 157306 710042 157542 710278
rect 153266 708442 153502 708678
rect 153586 708442 153822 708678
rect 153266 708122 153502 708358
rect 153586 708122 153822 708358
rect 149546 706522 149782 706758
rect 149866 706522 150102 706758
rect 149546 706202 149782 706438
rect 149866 706202 150102 706438
rect 138986 680378 139222 680614
rect 139306 680378 139542 680614
rect 138986 680058 139222 680294
rect 139306 680058 139542 680294
rect 138986 644378 139222 644614
rect 139306 644378 139542 644614
rect 138986 644058 139222 644294
rect 139306 644058 139542 644294
rect 138986 608378 139222 608614
rect 139306 608378 139542 608614
rect 138986 608058 139222 608294
rect 139306 608058 139542 608294
rect 138986 572378 139222 572614
rect 139306 572378 139542 572614
rect 138986 572058 139222 572294
rect 139306 572058 139542 572294
rect 138986 536378 139222 536614
rect 139306 536378 139542 536614
rect 138986 536058 139222 536294
rect 139306 536058 139542 536294
rect 138986 500378 139222 500614
rect 139306 500378 139542 500614
rect 138986 500058 139222 500294
rect 139306 500058 139542 500294
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 149546 654938 149782 655174
rect 149866 654938 150102 655174
rect 149546 654618 149782 654854
rect 149866 654618 150102 654854
rect 149546 618938 149782 619174
rect 149866 618938 150102 619174
rect 149546 618618 149782 618854
rect 149866 618618 150102 618854
rect 149546 582938 149782 583174
rect 149866 582938 150102 583174
rect 149546 582618 149782 582854
rect 149866 582618 150102 582854
rect 149546 546938 149782 547174
rect 149866 546938 150102 547174
rect 149546 546618 149782 546854
rect 149866 546618 150102 546854
rect 149546 510938 149782 511174
rect 149866 510938 150102 511174
rect 149546 510618 149782 510854
rect 149866 510618 150102 510854
rect 149546 474938 149782 475174
rect 149866 474938 150102 475174
rect 149546 474618 149782 474854
rect 149866 474618 150102 474854
rect 153266 694658 153502 694894
rect 153586 694658 153822 694894
rect 153266 694338 153502 694574
rect 153586 694338 153822 694574
rect 153266 658658 153502 658894
rect 153586 658658 153822 658894
rect 153266 658338 153502 658574
rect 153586 658338 153822 658574
rect 153266 622658 153502 622894
rect 153586 622658 153822 622894
rect 153266 622338 153502 622574
rect 153586 622338 153822 622574
rect 153266 586658 153502 586894
rect 153586 586658 153822 586894
rect 153266 586338 153502 586574
rect 153586 586338 153822 586574
rect 153266 550658 153502 550894
rect 153586 550658 153822 550894
rect 153266 550338 153502 550574
rect 153586 550338 153822 550574
rect 153266 514658 153502 514894
rect 153586 514658 153822 514894
rect 153266 514338 153502 514574
rect 153586 514338 153822 514574
rect 153266 478658 153502 478894
rect 153586 478658 153822 478894
rect 153266 478338 153502 478574
rect 153586 478338 153822 478574
rect 174986 711322 175222 711558
rect 175306 711322 175542 711558
rect 174986 711002 175222 711238
rect 175306 711002 175542 711238
rect 171266 709402 171502 709638
rect 171586 709402 171822 709638
rect 171266 709082 171502 709318
rect 171586 709082 171822 709318
rect 167546 707482 167782 707718
rect 167866 707482 168102 707718
rect 167546 707162 167782 707398
rect 167866 707162 168102 707398
rect 156986 698378 157222 698614
rect 157306 698378 157542 698614
rect 156986 698058 157222 698294
rect 157306 698058 157542 698294
rect 156986 662378 157222 662614
rect 157306 662378 157542 662614
rect 156986 662058 157222 662294
rect 157306 662058 157542 662294
rect 156986 626378 157222 626614
rect 157306 626378 157542 626614
rect 156986 626058 157222 626294
rect 157306 626058 157542 626294
rect 156986 590378 157222 590614
rect 157306 590378 157542 590614
rect 156986 590058 157222 590294
rect 157306 590058 157542 590294
rect 156986 554378 157222 554614
rect 157306 554378 157542 554614
rect 156986 554058 157222 554294
rect 157306 554058 157542 554294
rect 156986 518378 157222 518614
rect 157306 518378 157542 518614
rect 156986 518058 157222 518294
rect 157306 518058 157542 518294
rect 156986 482378 157222 482614
rect 157306 482378 157542 482614
rect 156986 482058 157222 482294
rect 157306 482058 157542 482294
rect 163826 705562 164062 705798
rect 164146 705562 164382 705798
rect 163826 705242 164062 705478
rect 164146 705242 164382 705478
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 163826 561218 164062 561454
rect 164146 561218 164382 561454
rect 163826 560898 164062 561134
rect 164146 560898 164382 561134
rect 163826 525218 164062 525454
rect 164146 525218 164382 525454
rect 163826 524898 164062 525134
rect 164146 524898 164382 525134
rect 163826 489218 164062 489454
rect 164146 489218 164382 489454
rect 163826 488898 164062 489134
rect 164146 488898 164382 489134
rect 167546 672938 167782 673174
rect 167866 672938 168102 673174
rect 167546 672618 167782 672854
rect 167866 672618 168102 672854
rect 167546 636938 167782 637174
rect 167866 636938 168102 637174
rect 167546 636618 167782 636854
rect 167866 636618 168102 636854
rect 167546 600938 167782 601174
rect 167866 600938 168102 601174
rect 167546 600618 167782 600854
rect 167866 600618 168102 600854
rect 167546 564938 167782 565174
rect 167866 564938 168102 565174
rect 167546 564618 167782 564854
rect 167866 564618 168102 564854
rect 167546 528938 167782 529174
rect 167866 528938 168102 529174
rect 167546 528618 167782 528854
rect 167866 528618 168102 528854
rect 167546 492938 167782 493174
rect 167866 492938 168102 493174
rect 167546 492618 167782 492854
rect 167866 492618 168102 492854
rect 171266 676658 171502 676894
rect 171586 676658 171822 676894
rect 171266 676338 171502 676574
rect 171586 676338 171822 676574
rect 171266 640658 171502 640894
rect 171586 640658 171822 640894
rect 171266 640338 171502 640574
rect 171586 640338 171822 640574
rect 171266 604658 171502 604894
rect 171586 604658 171822 604894
rect 171266 604338 171502 604574
rect 171586 604338 171822 604574
rect 171266 568658 171502 568894
rect 171586 568658 171822 568894
rect 171266 568338 171502 568574
rect 171586 568338 171822 568574
rect 171266 532658 171502 532894
rect 171586 532658 171822 532894
rect 171266 532338 171502 532574
rect 171586 532338 171822 532574
rect 171266 496658 171502 496894
rect 171586 496658 171822 496894
rect 171266 496338 171502 496574
rect 171586 496338 171822 496574
rect 192986 710362 193222 710598
rect 193306 710362 193542 710598
rect 192986 710042 193222 710278
rect 193306 710042 193542 710278
rect 189266 708442 189502 708678
rect 189586 708442 189822 708678
rect 189266 708122 189502 708358
rect 189586 708122 189822 708358
rect 185546 706522 185782 706758
rect 185866 706522 186102 706758
rect 185546 706202 185782 706438
rect 185866 706202 186102 706438
rect 174986 680378 175222 680614
rect 175306 680378 175542 680614
rect 174986 680058 175222 680294
rect 175306 680058 175542 680294
rect 174986 644378 175222 644614
rect 175306 644378 175542 644614
rect 174986 644058 175222 644294
rect 175306 644058 175542 644294
rect 174986 608378 175222 608614
rect 175306 608378 175542 608614
rect 174986 608058 175222 608294
rect 175306 608058 175542 608294
rect 174986 572378 175222 572614
rect 175306 572378 175542 572614
rect 174986 572058 175222 572294
rect 175306 572058 175542 572294
rect 174986 536378 175222 536614
rect 175306 536378 175542 536614
rect 174986 536058 175222 536294
rect 175306 536058 175542 536294
rect 174986 500378 175222 500614
rect 175306 500378 175542 500614
rect 174986 500058 175222 500294
rect 175306 500058 175542 500294
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 185546 690938 185782 691174
rect 185866 690938 186102 691174
rect 185546 690618 185782 690854
rect 185866 690618 186102 690854
rect 185546 654938 185782 655174
rect 185866 654938 186102 655174
rect 185546 654618 185782 654854
rect 185866 654618 186102 654854
rect 185546 618938 185782 619174
rect 185866 618938 186102 619174
rect 185546 618618 185782 618854
rect 185866 618618 186102 618854
rect 185546 582938 185782 583174
rect 185866 582938 186102 583174
rect 185546 582618 185782 582854
rect 185866 582618 186102 582854
rect 185546 546938 185782 547174
rect 185866 546938 186102 547174
rect 185546 546618 185782 546854
rect 185866 546618 186102 546854
rect 185546 510938 185782 511174
rect 185866 510938 186102 511174
rect 185546 510618 185782 510854
rect 185866 510618 186102 510854
rect 185546 474938 185782 475174
rect 185866 474938 186102 475174
rect 185546 474618 185782 474854
rect 185866 474618 186102 474854
rect 189266 694658 189502 694894
rect 189586 694658 189822 694894
rect 189266 694338 189502 694574
rect 189586 694338 189822 694574
rect 189266 658658 189502 658894
rect 189586 658658 189822 658894
rect 189266 658338 189502 658574
rect 189586 658338 189822 658574
rect 189266 622658 189502 622894
rect 189586 622658 189822 622894
rect 189266 622338 189502 622574
rect 189586 622338 189822 622574
rect 189266 586658 189502 586894
rect 189586 586658 189822 586894
rect 189266 586338 189502 586574
rect 189586 586338 189822 586574
rect 189266 550658 189502 550894
rect 189586 550658 189822 550894
rect 189266 550338 189502 550574
rect 189586 550338 189822 550574
rect 189266 514658 189502 514894
rect 189586 514658 189822 514894
rect 189266 514338 189502 514574
rect 189586 514338 189822 514574
rect 189266 478658 189502 478894
rect 189586 478658 189822 478894
rect 189266 478338 189502 478574
rect 189586 478338 189822 478574
rect 50328 453218 50564 453454
rect 50328 452898 50564 453134
rect 186056 453218 186292 453454
rect 186056 452898 186292 453134
rect 45266 442658 45502 442894
rect 45586 442658 45822 442894
rect 45266 442338 45502 442574
rect 45586 442338 45822 442574
rect 51008 435218 51244 435454
rect 51008 434898 51244 435134
rect 185376 435218 185612 435454
rect 185376 434898 185612 435134
rect 50328 417218 50564 417454
rect 50328 416898 50564 417134
rect 186056 417218 186292 417454
rect 186056 416898 186292 417134
rect 45266 406658 45502 406894
rect 45586 406658 45822 406894
rect 45266 406338 45502 406574
rect 45586 406338 45822 406574
rect 51008 399218 51244 399454
rect 51008 398898 51244 399134
rect 185376 399218 185612 399454
rect 185376 398898 185612 399134
rect 50328 381218 50564 381454
rect 50328 380898 50564 381134
rect 186056 381218 186292 381454
rect 186056 380898 186292 381134
rect 45266 370658 45502 370894
rect 45586 370658 45822 370894
rect 45266 370338 45502 370574
rect 45586 370338 45822 370574
rect 45266 334658 45502 334894
rect 45586 334658 45822 334894
rect 45266 334338 45502 334574
rect 45586 334338 45822 334574
rect 45266 298658 45502 298894
rect 45586 298658 45822 298894
rect 45266 298338 45502 298574
rect 45586 298338 45822 298574
rect 48986 374378 49222 374614
rect 49306 374378 49542 374614
rect 48986 374058 49222 374294
rect 49306 374058 49542 374294
rect 48986 338378 49222 338614
rect 49306 338378 49542 338614
rect 48986 338058 49222 338294
rect 49306 338058 49542 338294
rect 48986 302378 49222 302614
rect 49306 302378 49542 302614
rect 48986 302058 49222 302294
rect 49306 302058 49542 302294
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 59546 348938 59782 349174
rect 59866 348938 60102 349174
rect 59546 348618 59782 348854
rect 59866 348618 60102 348854
rect 59546 312938 59782 313174
rect 59866 312938 60102 313174
rect 59546 312618 59782 312854
rect 59866 312618 60102 312854
rect 63266 352658 63502 352894
rect 63586 352658 63822 352894
rect 63266 352338 63502 352574
rect 63586 352338 63822 352574
rect 63266 316658 63502 316894
rect 63586 316658 63822 316894
rect 63266 316338 63502 316574
rect 63586 316338 63822 316574
rect 66986 356378 67222 356614
rect 67306 356378 67542 356614
rect 66986 356058 67222 356294
rect 67306 356058 67542 356294
rect 66986 320378 67222 320614
rect 67306 320378 67542 320614
rect 66986 320058 67222 320294
rect 67306 320058 67542 320294
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 73826 327218 74062 327454
rect 74146 327218 74382 327454
rect 73826 326898 74062 327134
rect 74146 326898 74382 327134
rect 73826 291218 74062 291454
rect 74146 291218 74382 291454
rect 73826 290898 74062 291134
rect 74146 290898 74382 291134
rect 77546 366938 77782 367174
rect 77866 366938 78102 367174
rect 77546 366618 77782 366854
rect 77866 366618 78102 366854
rect 77546 330938 77782 331174
rect 77866 330938 78102 331174
rect 77546 330618 77782 330854
rect 77866 330618 78102 330854
rect 77546 294938 77782 295174
rect 77866 294938 78102 295174
rect 77546 294618 77782 294854
rect 77866 294618 78102 294854
rect 81266 370658 81502 370894
rect 81586 370658 81822 370894
rect 81266 370338 81502 370574
rect 81586 370338 81822 370574
rect 81266 334658 81502 334894
rect 81586 334658 81822 334894
rect 81266 334338 81502 334574
rect 81586 334338 81822 334574
rect 81266 298658 81502 298894
rect 81586 298658 81822 298894
rect 81266 298338 81502 298574
rect 81586 298338 81822 298574
rect 84986 374378 85222 374614
rect 85306 374378 85542 374614
rect 84986 374058 85222 374294
rect 85306 374058 85542 374294
rect 84986 338378 85222 338614
rect 85306 338378 85542 338614
rect 84986 338058 85222 338294
rect 85306 338058 85542 338294
rect 84986 302378 85222 302614
rect 85306 302378 85542 302614
rect 84986 302058 85222 302294
rect 85306 302058 85542 302294
rect 91826 345218 92062 345454
rect 92146 345218 92382 345454
rect 91826 344898 92062 345134
rect 92146 344898 92382 345134
rect 91826 309218 92062 309454
rect 92146 309218 92382 309454
rect 91826 308898 92062 309134
rect 92146 308898 92382 309134
rect 95546 348938 95782 349174
rect 95866 348938 96102 349174
rect 95546 348618 95782 348854
rect 95866 348618 96102 348854
rect 95546 312938 95782 313174
rect 95866 312938 96102 313174
rect 95546 312618 95782 312854
rect 95866 312618 96102 312854
rect 99266 352658 99502 352894
rect 99586 352658 99822 352894
rect 99266 352338 99502 352574
rect 99586 352338 99822 352574
rect 99266 316658 99502 316894
rect 99586 316658 99822 316894
rect 99266 316338 99502 316574
rect 99586 316338 99822 316574
rect 102986 356378 103222 356614
rect 103306 356378 103542 356614
rect 102986 356058 103222 356294
rect 103306 356058 103542 356294
rect 102986 320378 103222 320614
rect 103306 320378 103542 320614
rect 102986 320058 103222 320294
rect 103306 320058 103542 320294
rect 109826 363218 110062 363454
rect 110146 363218 110382 363454
rect 109826 362898 110062 363134
rect 110146 362898 110382 363134
rect 109826 327218 110062 327454
rect 110146 327218 110382 327454
rect 109826 326898 110062 327134
rect 110146 326898 110382 327134
rect 109826 291218 110062 291454
rect 110146 291218 110382 291454
rect 109826 290898 110062 291134
rect 110146 290898 110382 291134
rect 113546 366938 113782 367174
rect 113866 366938 114102 367174
rect 113546 366618 113782 366854
rect 113866 366618 114102 366854
rect 113546 330938 113782 331174
rect 113866 330938 114102 331174
rect 113546 330618 113782 330854
rect 113866 330618 114102 330854
rect 113546 294938 113782 295174
rect 113866 294938 114102 295174
rect 113546 294618 113782 294854
rect 113866 294618 114102 294854
rect 117266 370658 117502 370894
rect 117586 370658 117822 370894
rect 117266 370338 117502 370574
rect 117586 370338 117822 370574
rect 117266 334658 117502 334894
rect 117586 334658 117822 334894
rect 117266 334338 117502 334574
rect 117586 334338 117822 334574
rect 117266 298658 117502 298894
rect 117586 298658 117822 298894
rect 117266 298338 117502 298574
rect 117586 298338 117822 298574
rect 120986 374378 121222 374614
rect 121306 374378 121542 374614
rect 120986 374058 121222 374294
rect 121306 374058 121542 374294
rect 120986 338378 121222 338614
rect 121306 338378 121542 338614
rect 120986 338058 121222 338294
rect 121306 338058 121542 338294
rect 120986 302378 121222 302614
rect 121306 302378 121542 302614
rect 120986 302058 121222 302294
rect 121306 302058 121542 302294
rect 127826 345218 128062 345454
rect 128146 345218 128382 345454
rect 127826 344898 128062 345134
rect 128146 344898 128382 345134
rect 127826 309218 128062 309454
rect 128146 309218 128382 309454
rect 127826 308898 128062 309134
rect 128146 308898 128382 309134
rect 131546 348938 131782 349174
rect 131866 348938 132102 349174
rect 131546 348618 131782 348854
rect 131866 348618 132102 348854
rect 131546 312938 131782 313174
rect 131866 312938 132102 313174
rect 131546 312618 131782 312854
rect 131866 312618 132102 312854
rect 135266 352658 135502 352894
rect 135586 352658 135822 352894
rect 135266 352338 135502 352574
rect 135586 352338 135822 352574
rect 135266 316658 135502 316894
rect 135586 316658 135822 316894
rect 135266 316338 135502 316574
rect 135586 316338 135822 316574
rect 138986 356378 139222 356614
rect 139306 356378 139542 356614
rect 138986 356058 139222 356294
rect 139306 356058 139542 356294
rect 138986 320378 139222 320614
rect 139306 320378 139542 320614
rect 138986 320058 139222 320294
rect 139306 320058 139542 320294
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 145826 327218 146062 327454
rect 146146 327218 146382 327454
rect 145826 326898 146062 327134
rect 146146 326898 146382 327134
rect 145826 291218 146062 291454
rect 146146 291218 146382 291454
rect 145826 290898 146062 291134
rect 146146 290898 146382 291134
rect 149546 366938 149782 367174
rect 149866 366938 150102 367174
rect 149546 366618 149782 366854
rect 149866 366618 150102 366854
rect 149546 330938 149782 331174
rect 149866 330938 150102 331174
rect 149546 330618 149782 330854
rect 149866 330618 150102 330854
rect 149546 294938 149782 295174
rect 149866 294938 150102 295174
rect 149546 294618 149782 294854
rect 149866 294618 150102 294854
rect 153266 370658 153502 370894
rect 153586 370658 153822 370894
rect 153266 370338 153502 370574
rect 153586 370338 153822 370574
rect 153266 334658 153502 334894
rect 153586 334658 153822 334894
rect 153266 334338 153502 334574
rect 153586 334338 153822 334574
rect 153266 298658 153502 298894
rect 153586 298658 153822 298894
rect 153266 298338 153502 298574
rect 153586 298338 153822 298574
rect 156986 374378 157222 374614
rect 157306 374378 157542 374614
rect 156986 374058 157222 374294
rect 157306 374058 157542 374294
rect 156986 338378 157222 338614
rect 157306 338378 157542 338614
rect 156986 338058 157222 338294
rect 157306 338058 157542 338294
rect 156986 302378 157222 302614
rect 157306 302378 157542 302614
rect 156986 302058 157222 302294
rect 157306 302058 157542 302294
rect 163826 345218 164062 345454
rect 164146 345218 164382 345454
rect 163826 344898 164062 345134
rect 164146 344898 164382 345134
rect 163826 309218 164062 309454
rect 164146 309218 164382 309454
rect 163826 308898 164062 309134
rect 164146 308898 164382 309134
rect 167546 348938 167782 349174
rect 167866 348938 168102 349174
rect 167546 348618 167782 348854
rect 167866 348618 168102 348854
rect 167546 312938 167782 313174
rect 167866 312938 168102 313174
rect 167546 312618 167782 312854
rect 167866 312618 168102 312854
rect 171266 352658 171502 352894
rect 171586 352658 171822 352894
rect 171266 352338 171502 352574
rect 171586 352338 171822 352574
rect 171266 316658 171502 316894
rect 171586 316658 171822 316894
rect 171266 316338 171502 316574
rect 171586 316338 171822 316574
rect 174986 356378 175222 356614
rect 175306 356378 175542 356614
rect 174986 356058 175222 356294
rect 175306 356058 175542 356294
rect 174986 320378 175222 320614
rect 175306 320378 175542 320614
rect 174986 320058 175222 320294
rect 175306 320058 175542 320294
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 181826 327218 182062 327454
rect 182146 327218 182382 327454
rect 181826 326898 182062 327134
rect 182146 326898 182382 327134
rect 181826 291218 182062 291454
rect 182146 291218 182382 291454
rect 181826 290898 182062 291134
rect 182146 290898 182382 291134
rect 185546 366938 185782 367174
rect 185866 366938 186102 367174
rect 185546 366618 185782 366854
rect 185866 366618 186102 366854
rect 185546 330938 185782 331174
rect 185866 330938 186102 331174
rect 185546 330618 185782 330854
rect 185866 330618 186102 330854
rect 189266 442658 189502 442894
rect 189586 442658 189822 442894
rect 189266 442338 189502 442574
rect 189586 442338 189822 442574
rect 189266 406658 189502 406894
rect 189586 406658 189822 406894
rect 189266 406338 189502 406574
rect 189586 406338 189822 406574
rect 189266 370658 189502 370894
rect 189586 370658 189822 370894
rect 189266 370338 189502 370574
rect 189586 370338 189822 370574
rect 189266 334658 189502 334894
rect 189586 334658 189822 334894
rect 189266 334338 189502 334574
rect 189586 334338 189822 334574
rect 185546 294938 185782 295174
rect 185866 294938 186102 295174
rect 185546 294618 185782 294854
rect 185866 294618 186102 294854
rect 189266 298658 189502 298894
rect 189586 298658 189822 298894
rect 189266 298338 189502 298574
rect 189586 298338 189822 298574
rect 50328 273218 50564 273454
rect 50328 272898 50564 273134
rect 186056 273218 186292 273454
rect 186056 272898 186292 273134
rect 45266 262658 45502 262894
rect 45586 262658 45822 262894
rect 45266 262338 45502 262574
rect 45586 262338 45822 262574
rect 51008 255218 51244 255454
rect 51008 254898 51244 255134
rect 185376 255218 185612 255454
rect 185376 254898 185612 255134
rect 50328 237218 50564 237454
rect 50328 236898 50564 237134
rect 186056 237218 186292 237454
rect 186056 236898 186292 237134
rect 45266 226658 45502 226894
rect 45586 226658 45822 226894
rect 45266 226338 45502 226574
rect 45586 226338 45822 226574
rect 51008 219218 51244 219454
rect 51008 218898 51244 219134
rect 185376 219218 185612 219454
rect 185376 218898 185612 219134
rect 50328 201218 50564 201454
rect 50328 200898 50564 201134
rect 186056 201218 186292 201454
rect 186056 200898 186292 201134
rect 45266 190658 45502 190894
rect 45586 190658 45822 190894
rect 45266 190338 45502 190574
rect 45586 190338 45822 190574
rect 45266 154658 45502 154894
rect 45586 154658 45822 154894
rect 45266 154338 45502 154574
rect 45586 154338 45822 154574
rect 45266 118658 45502 118894
rect 45586 118658 45822 118894
rect 45266 118338 45502 118574
rect 45586 118338 45822 118574
rect 45266 82658 45502 82894
rect 45586 82658 45822 82894
rect 45266 82338 45502 82574
rect 45586 82338 45822 82574
rect 45266 46658 45502 46894
rect 45586 46658 45822 46894
rect 45266 46338 45502 46574
rect 45586 46338 45822 46574
rect 45266 10658 45502 10894
rect 45586 10658 45822 10894
rect 45266 10338 45502 10574
rect 45586 10338 45822 10574
rect 45266 -4422 45502 -4186
rect 45586 -4422 45822 -4186
rect 45266 -4742 45502 -4506
rect 45586 -4742 45822 -4506
rect 48986 194378 49222 194614
rect 49306 194378 49542 194614
rect 48986 194058 49222 194294
rect 49306 194058 49542 194294
rect 48986 158378 49222 158614
rect 49306 158378 49542 158614
rect 48986 158058 49222 158294
rect 49306 158058 49542 158294
rect 48986 122378 49222 122614
rect 49306 122378 49542 122614
rect 48986 122058 49222 122294
rect 49306 122058 49542 122294
rect 48986 86378 49222 86614
rect 49306 86378 49542 86614
rect 48986 86058 49222 86294
rect 49306 86058 49542 86294
rect 48986 50378 49222 50614
rect 49306 50378 49542 50614
rect 48986 50058 49222 50294
rect 49306 50058 49542 50294
rect 48986 14378 49222 14614
rect 49306 14378 49542 14614
rect 48986 14058 49222 14294
rect 49306 14058 49542 14294
rect 30986 -7302 31222 -7066
rect 31306 -7302 31542 -7066
rect 30986 -7622 31222 -7386
rect 31306 -7622 31542 -7386
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -1542 56062 -1306
rect 56146 -1542 56382 -1306
rect 55826 -1862 56062 -1626
rect 56146 -1862 56382 -1626
rect 59546 168938 59782 169174
rect 59866 168938 60102 169174
rect 59546 168618 59782 168854
rect 59866 168618 60102 168854
rect 59546 132938 59782 133174
rect 59866 132938 60102 133174
rect 59546 132618 59782 132854
rect 59866 132618 60102 132854
rect 59546 96938 59782 97174
rect 59866 96938 60102 97174
rect 59546 96618 59782 96854
rect 59866 96618 60102 96854
rect 59546 60938 59782 61174
rect 59866 60938 60102 61174
rect 59546 60618 59782 60854
rect 59866 60618 60102 60854
rect 59546 24938 59782 25174
rect 59866 24938 60102 25174
rect 59546 24618 59782 24854
rect 59866 24618 60102 24854
rect 59546 -3462 59782 -3226
rect 59866 -3462 60102 -3226
rect 59546 -3782 59782 -3546
rect 59866 -3782 60102 -3546
rect 63266 172658 63502 172894
rect 63586 172658 63822 172894
rect 63266 172338 63502 172574
rect 63586 172338 63822 172574
rect 63266 136658 63502 136894
rect 63586 136658 63822 136894
rect 63266 136338 63502 136574
rect 63586 136338 63822 136574
rect 63266 100658 63502 100894
rect 63586 100658 63822 100894
rect 63266 100338 63502 100574
rect 63586 100338 63822 100574
rect 63266 64658 63502 64894
rect 63586 64658 63822 64894
rect 63266 64338 63502 64574
rect 63586 64338 63822 64574
rect 63266 28658 63502 28894
rect 63586 28658 63822 28894
rect 63266 28338 63502 28574
rect 63586 28338 63822 28574
rect 63266 -5382 63502 -5146
rect 63586 -5382 63822 -5146
rect 63266 -5702 63502 -5466
rect 63586 -5702 63822 -5466
rect 66986 176378 67222 176614
rect 67306 176378 67542 176614
rect 66986 176058 67222 176294
rect 67306 176058 67542 176294
rect 66986 140378 67222 140614
rect 67306 140378 67542 140614
rect 66986 140058 67222 140294
rect 67306 140058 67542 140294
rect 66986 104378 67222 104614
rect 67306 104378 67542 104614
rect 66986 104058 67222 104294
rect 67306 104058 67542 104294
rect 66986 68378 67222 68614
rect 67306 68378 67542 68614
rect 66986 68058 67222 68294
rect 67306 68058 67542 68294
rect 66986 32378 67222 32614
rect 67306 32378 67542 32614
rect 66986 32058 67222 32294
rect 67306 32058 67542 32294
rect 48986 -6342 49222 -6106
rect 49306 -6342 49542 -6106
rect 48986 -6662 49222 -6426
rect 49306 -6662 49542 -6426
rect 73826 183218 74062 183454
rect 74146 183218 74382 183454
rect 73826 182898 74062 183134
rect 74146 182898 74382 183134
rect 73826 147218 74062 147454
rect 74146 147218 74382 147454
rect 73826 146898 74062 147134
rect 74146 146898 74382 147134
rect 73826 111218 74062 111454
rect 74146 111218 74382 111454
rect 73826 110898 74062 111134
rect 74146 110898 74382 111134
rect 73826 75218 74062 75454
rect 74146 75218 74382 75454
rect 73826 74898 74062 75134
rect 74146 74898 74382 75134
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 186938 77782 187174
rect 77866 186938 78102 187174
rect 77546 186618 77782 186854
rect 77866 186618 78102 186854
rect 77546 150938 77782 151174
rect 77866 150938 78102 151174
rect 77546 150618 77782 150854
rect 77866 150618 78102 150854
rect 77546 114938 77782 115174
rect 77866 114938 78102 115174
rect 77546 114618 77782 114854
rect 77866 114618 78102 114854
rect 77546 78938 77782 79174
rect 77866 78938 78102 79174
rect 77546 78618 77782 78854
rect 77866 78618 78102 78854
rect 77546 42938 77782 43174
rect 77866 42938 78102 43174
rect 77546 42618 77782 42854
rect 77866 42618 78102 42854
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -2502 77782 -2266
rect 77866 -2502 78102 -2266
rect 77546 -2822 77782 -2586
rect 77866 -2822 78102 -2586
rect 81266 190658 81502 190894
rect 81586 190658 81822 190894
rect 81266 190338 81502 190574
rect 81586 190338 81822 190574
rect 81266 154658 81502 154894
rect 81586 154658 81822 154894
rect 81266 154338 81502 154574
rect 81586 154338 81822 154574
rect 81266 118658 81502 118894
rect 81586 118658 81822 118894
rect 81266 118338 81502 118574
rect 81586 118338 81822 118574
rect 81266 82658 81502 82894
rect 81586 82658 81822 82894
rect 81266 82338 81502 82574
rect 81586 82338 81822 82574
rect 81266 46658 81502 46894
rect 81586 46658 81822 46894
rect 81266 46338 81502 46574
rect 81586 46338 81822 46574
rect 81266 10658 81502 10894
rect 81586 10658 81822 10894
rect 81266 10338 81502 10574
rect 81586 10338 81822 10574
rect 81266 -4422 81502 -4186
rect 81586 -4422 81822 -4186
rect 81266 -4742 81502 -4506
rect 81586 -4742 81822 -4506
rect 84986 194378 85222 194614
rect 85306 194378 85542 194614
rect 84986 194058 85222 194294
rect 85306 194058 85542 194294
rect 84986 158378 85222 158614
rect 85306 158378 85542 158614
rect 84986 158058 85222 158294
rect 85306 158058 85542 158294
rect 84986 122378 85222 122614
rect 85306 122378 85542 122614
rect 84986 122058 85222 122294
rect 85306 122058 85542 122294
rect 84986 86378 85222 86614
rect 85306 86378 85542 86614
rect 84986 86058 85222 86294
rect 85306 86058 85542 86294
rect 84986 50378 85222 50614
rect 85306 50378 85542 50614
rect 84986 50058 85222 50294
rect 85306 50058 85542 50294
rect 84986 14378 85222 14614
rect 85306 14378 85542 14614
rect 84986 14058 85222 14294
rect 85306 14058 85542 14294
rect 66986 -7302 67222 -7066
rect 67306 -7302 67542 -7066
rect 66986 -7622 67222 -7386
rect 67306 -7622 67542 -7386
rect 91826 165218 92062 165454
rect 92146 165218 92382 165454
rect 91826 164898 92062 165134
rect 92146 164898 92382 165134
rect 91826 129218 92062 129454
rect 92146 129218 92382 129454
rect 91826 128898 92062 129134
rect 92146 128898 92382 129134
rect 91826 93218 92062 93454
rect 92146 93218 92382 93454
rect 91826 92898 92062 93134
rect 92146 92898 92382 93134
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -1542 92062 -1306
rect 92146 -1542 92382 -1306
rect 91826 -1862 92062 -1626
rect 92146 -1862 92382 -1626
rect 95546 168938 95782 169174
rect 95866 168938 96102 169174
rect 95546 168618 95782 168854
rect 95866 168618 96102 168854
rect 95546 132938 95782 133174
rect 95866 132938 96102 133174
rect 95546 132618 95782 132854
rect 95866 132618 96102 132854
rect 95546 96938 95782 97174
rect 95866 96938 96102 97174
rect 95546 96618 95782 96854
rect 95866 96618 96102 96854
rect 95546 60938 95782 61174
rect 95866 60938 96102 61174
rect 95546 60618 95782 60854
rect 95866 60618 96102 60854
rect 95546 24938 95782 25174
rect 95866 24938 96102 25174
rect 95546 24618 95782 24854
rect 95866 24618 96102 24854
rect 95546 -3462 95782 -3226
rect 95866 -3462 96102 -3226
rect 95546 -3782 95782 -3546
rect 95866 -3782 96102 -3546
rect 99266 172658 99502 172894
rect 99586 172658 99822 172894
rect 99266 172338 99502 172574
rect 99586 172338 99822 172574
rect 99266 136658 99502 136894
rect 99586 136658 99822 136894
rect 99266 136338 99502 136574
rect 99586 136338 99822 136574
rect 99266 100658 99502 100894
rect 99586 100658 99822 100894
rect 99266 100338 99502 100574
rect 99586 100338 99822 100574
rect 99266 64658 99502 64894
rect 99586 64658 99822 64894
rect 99266 64338 99502 64574
rect 99586 64338 99822 64574
rect 99266 28658 99502 28894
rect 99586 28658 99822 28894
rect 99266 28338 99502 28574
rect 99586 28338 99822 28574
rect 99266 -5382 99502 -5146
rect 99586 -5382 99822 -5146
rect 99266 -5702 99502 -5466
rect 99586 -5702 99822 -5466
rect 102986 176378 103222 176614
rect 103306 176378 103542 176614
rect 102986 176058 103222 176294
rect 103306 176058 103542 176294
rect 102986 140378 103222 140614
rect 103306 140378 103542 140614
rect 102986 140058 103222 140294
rect 103306 140058 103542 140294
rect 102986 104378 103222 104614
rect 103306 104378 103542 104614
rect 102986 104058 103222 104294
rect 103306 104058 103542 104294
rect 102986 68378 103222 68614
rect 103306 68378 103542 68614
rect 102986 68058 103222 68294
rect 103306 68058 103542 68294
rect 102986 32378 103222 32614
rect 103306 32378 103542 32614
rect 102986 32058 103222 32294
rect 103306 32058 103542 32294
rect 84986 -6342 85222 -6106
rect 85306 -6342 85542 -6106
rect 84986 -6662 85222 -6426
rect 85306 -6662 85542 -6426
rect 109826 183218 110062 183454
rect 110146 183218 110382 183454
rect 109826 182898 110062 183134
rect 110146 182898 110382 183134
rect 109826 147218 110062 147454
rect 110146 147218 110382 147454
rect 109826 146898 110062 147134
rect 110146 146898 110382 147134
rect 109826 111218 110062 111454
rect 110146 111218 110382 111454
rect 109826 110898 110062 111134
rect 110146 110898 110382 111134
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 186938 113782 187174
rect 113866 186938 114102 187174
rect 113546 186618 113782 186854
rect 113866 186618 114102 186854
rect 113546 150938 113782 151174
rect 113866 150938 114102 151174
rect 113546 150618 113782 150854
rect 113866 150618 114102 150854
rect 113546 114938 113782 115174
rect 113866 114938 114102 115174
rect 113546 114618 113782 114854
rect 113866 114618 114102 114854
rect 113546 78938 113782 79174
rect 113866 78938 114102 79174
rect 113546 78618 113782 78854
rect 113866 78618 114102 78854
rect 113546 42938 113782 43174
rect 113866 42938 114102 43174
rect 113546 42618 113782 42854
rect 113866 42618 114102 42854
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 113546 -2502 113782 -2266
rect 113866 -2502 114102 -2266
rect 113546 -2822 113782 -2586
rect 113866 -2822 114102 -2586
rect 117266 190658 117502 190894
rect 117586 190658 117822 190894
rect 117266 190338 117502 190574
rect 117586 190338 117822 190574
rect 117266 154658 117502 154894
rect 117586 154658 117822 154894
rect 117266 154338 117502 154574
rect 117586 154338 117822 154574
rect 117266 118658 117502 118894
rect 117586 118658 117822 118894
rect 117266 118338 117502 118574
rect 117586 118338 117822 118574
rect 117266 82658 117502 82894
rect 117586 82658 117822 82894
rect 117266 82338 117502 82574
rect 117586 82338 117822 82574
rect 117266 46658 117502 46894
rect 117586 46658 117822 46894
rect 117266 46338 117502 46574
rect 117586 46338 117822 46574
rect 117266 10658 117502 10894
rect 117586 10658 117822 10894
rect 117266 10338 117502 10574
rect 117586 10338 117822 10574
rect 117266 -4422 117502 -4186
rect 117586 -4422 117822 -4186
rect 117266 -4742 117502 -4506
rect 117586 -4742 117822 -4506
rect 120986 194378 121222 194614
rect 121306 194378 121542 194614
rect 120986 194058 121222 194294
rect 121306 194058 121542 194294
rect 120986 158378 121222 158614
rect 121306 158378 121542 158614
rect 120986 158058 121222 158294
rect 121306 158058 121542 158294
rect 120986 122378 121222 122614
rect 121306 122378 121542 122614
rect 120986 122058 121222 122294
rect 121306 122058 121542 122294
rect 120986 86378 121222 86614
rect 121306 86378 121542 86614
rect 120986 86058 121222 86294
rect 121306 86058 121542 86294
rect 120986 50378 121222 50614
rect 121306 50378 121542 50614
rect 120986 50058 121222 50294
rect 121306 50058 121542 50294
rect 120986 14378 121222 14614
rect 121306 14378 121542 14614
rect 120986 14058 121222 14294
rect 121306 14058 121542 14294
rect 102986 -7302 103222 -7066
rect 103306 -7302 103542 -7066
rect 102986 -7622 103222 -7386
rect 103306 -7622 103542 -7386
rect 127826 165218 128062 165454
rect 128146 165218 128382 165454
rect 127826 164898 128062 165134
rect 128146 164898 128382 165134
rect 127826 129218 128062 129454
rect 128146 129218 128382 129454
rect 127826 128898 128062 129134
rect 128146 128898 128382 129134
rect 127826 93218 128062 93454
rect 128146 93218 128382 93454
rect 127826 92898 128062 93134
rect 128146 92898 128382 93134
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -1542 128062 -1306
rect 128146 -1542 128382 -1306
rect 127826 -1862 128062 -1626
rect 128146 -1862 128382 -1626
rect 131546 168938 131782 169174
rect 131866 168938 132102 169174
rect 131546 168618 131782 168854
rect 131866 168618 132102 168854
rect 131546 132938 131782 133174
rect 131866 132938 132102 133174
rect 131546 132618 131782 132854
rect 131866 132618 132102 132854
rect 131546 96938 131782 97174
rect 131866 96938 132102 97174
rect 131546 96618 131782 96854
rect 131866 96618 132102 96854
rect 131546 60938 131782 61174
rect 131866 60938 132102 61174
rect 131546 60618 131782 60854
rect 131866 60618 132102 60854
rect 131546 24938 131782 25174
rect 131866 24938 132102 25174
rect 131546 24618 131782 24854
rect 131866 24618 132102 24854
rect 131546 -3462 131782 -3226
rect 131866 -3462 132102 -3226
rect 131546 -3782 131782 -3546
rect 131866 -3782 132102 -3546
rect 135266 172658 135502 172894
rect 135586 172658 135822 172894
rect 135266 172338 135502 172574
rect 135586 172338 135822 172574
rect 135266 136658 135502 136894
rect 135586 136658 135822 136894
rect 135266 136338 135502 136574
rect 135586 136338 135822 136574
rect 135266 100658 135502 100894
rect 135586 100658 135822 100894
rect 135266 100338 135502 100574
rect 135586 100338 135822 100574
rect 135266 64658 135502 64894
rect 135586 64658 135822 64894
rect 135266 64338 135502 64574
rect 135586 64338 135822 64574
rect 135266 28658 135502 28894
rect 135586 28658 135822 28894
rect 135266 28338 135502 28574
rect 135586 28338 135822 28574
rect 135266 -5382 135502 -5146
rect 135586 -5382 135822 -5146
rect 135266 -5702 135502 -5466
rect 135586 -5702 135822 -5466
rect 138986 176378 139222 176614
rect 139306 176378 139542 176614
rect 138986 176058 139222 176294
rect 139306 176058 139542 176294
rect 138986 140378 139222 140614
rect 139306 140378 139542 140614
rect 138986 140058 139222 140294
rect 139306 140058 139542 140294
rect 138986 104378 139222 104614
rect 139306 104378 139542 104614
rect 138986 104058 139222 104294
rect 139306 104058 139542 104294
rect 138986 68378 139222 68614
rect 139306 68378 139542 68614
rect 138986 68058 139222 68294
rect 139306 68058 139542 68294
rect 138986 32378 139222 32614
rect 139306 32378 139542 32614
rect 138986 32058 139222 32294
rect 139306 32058 139542 32294
rect 120986 -6342 121222 -6106
rect 121306 -6342 121542 -6106
rect 120986 -6662 121222 -6426
rect 121306 -6662 121542 -6426
rect 145826 183218 146062 183454
rect 146146 183218 146382 183454
rect 145826 182898 146062 183134
rect 146146 182898 146382 183134
rect 145826 147218 146062 147454
rect 146146 147218 146382 147454
rect 145826 146898 146062 147134
rect 146146 146898 146382 147134
rect 145826 111218 146062 111454
rect 146146 111218 146382 111454
rect 145826 110898 146062 111134
rect 146146 110898 146382 111134
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 186938 149782 187174
rect 149866 186938 150102 187174
rect 149546 186618 149782 186854
rect 149866 186618 150102 186854
rect 149546 150938 149782 151174
rect 149866 150938 150102 151174
rect 149546 150618 149782 150854
rect 149866 150618 150102 150854
rect 149546 114938 149782 115174
rect 149866 114938 150102 115174
rect 149546 114618 149782 114854
rect 149866 114618 150102 114854
rect 149546 78938 149782 79174
rect 149866 78938 150102 79174
rect 149546 78618 149782 78854
rect 149866 78618 150102 78854
rect 149546 42938 149782 43174
rect 149866 42938 150102 43174
rect 149546 42618 149782 42854
rect 149866 42618 150102 42854
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 149546 -2502 149782 -2266
rect 149866 -2502 150102 -2266
rect 149546 -2822 149782 -2586
rect 149866 -2822 150102 -2586
rect 153266 190658 153502 190894
rect 153586 190658 153822 190894
rect 153266 190338 153502 190574
rect 153586 190338 153822 190574
rect 153266 154658 153502 154894
rect 153586 154658 153822 154894
rect 153266 154338 153502 154574
rect 153586 154338 153822 154574
rect 153266 118658 153502 118894
rect 153586 118658 153822 118894
rect 153266 118338 153502 118574
rect 153586 118338 153822 118574
rect 153266 82658 153502 82894
rect 153586 82658 153822 82894
rect 153266 82338 153502 82574
rect 153586 82338 153822 82574
rect 153266 46658 153502 46894
rect 153586 46658 153822 46894
rect 153266 46338 153502 46574
rect 153586 46338 153822 46574
rect 153266 10658 153502 10894
rect 153586 10658 153822 10894
rect 153266 10338 153502 10574
rect 153586 10338 153822 10574
rect 153266 -4422 153502 -4186
rect 153586 -4422 153822 -4186
rect 153266 -4742 153502 -4506
rect 153586 -4742 153822 -4506
rect 156986 194378 157222 194614
rect 157306 194378 157542 194614
rect 156986 194058 157222 194294
rect 157306 194058 157542 194294
rect 156986 158378 157222 158614
rect 157306 158378 157542 158614
rect 156986 158058 157222 158294
rect 157306 158058 157542 158294
rect 156986 122378 157222 122614
rect 157306 122378 157542 122614
rect 156986 122058 157222 122294
rect 157306 122058 157542 122294
rect 156986 86378 157222 86614
rect 157306 86378 157542 86614
rect 156986 86058 157222 86294
rect 157306 86058 157542 86294
rect 156986 50378 157222 50614
rect 157306 50378 157542 50614
rect 156986 50058 157222 50294
rect 157306 50058 157542 50294
rect 156986 14378 157222 14614
rect 157306 14378 157542 14614
rect 156986 14058 157222 14294
rect 157306 14058 157542 14294
rect 138986 -7302 139222 -7066
rect 139306 -7302 139542 -7066
rect 138986 -7622 139222 -7386
rect 139306 -7622 139542 -7386
rect 163826 165218 164062 165454
rect 164146 165218 164382 165454
rect 163826 164898 164062 165134
rect 164146 164898 164382 165134
rect 163826 129218 164062 129454
rect 164146 129218 164382 129454
rect 163826 128898 164062 129134
rect 164146 128898 164382 129134
rect 163826 93218 164062 93454
rect 164146 93218 164382 93454
rect 163826 92898 164062 93134
rect 164146 92898 164382 93134
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -1542 164062 -1306
rect 164146 -1542 164382 -1306
rect 163826 -1862 164062 -1626
rect 164146 -1862 164382 -1626
rect 167546 168938 167782 169174
rect 167866 168938 168102 169174
rect 167546 168618 167782 168854
rect 167866 168618 168102 168854
rect 167546 132938 167782 133174
rect 167866 132938 168102 133174
rect 167546 132618 167782 132854
rect 167866 132618 168102 132854
rect 167546 96938 167782 97174
rect 167866 96938 168102 97174
rect 167546 96618 167782 96854
rect 167866 96618 168102 96854
rect 167546 60938 167782 61174
rect 167866 60938 168102 61174
rect 167546 60618 167782 60854
rect 167866 60618 168102 60854
rect 167546 24938 167782 25174
rect 167866 24938 168102 25174
rect 167546 24618 167782 24854
rect 167866 24618 168102 24854
rect 167546 -3462 167782 -3226
rect 167866 -3462 168102 -3226
rect 167546 -3782 167782 -3546
rect 167866 -3782 168102 -3546
rect 189266 262658 189502 262894
rect 189586 262658 189822 262894
rect 189266 262338 189502 262574
rect 189586 262338 189822 262574
rect 189266 226658 189502 226894
rect 189586 226658 189822 226894
rect 189266 226338 189502 226574
rect 189586 226338 189822 226574
rect 171266 172658 171502 172894
rect 171586 172658 171822 172894
rect 171266 172338 171502 172574
rect 171586 172338 171822 172574
rect 171266 136658 171502 136894
rect 171586 136658 171822 136894
rect 171266 136338 171502 136574
rect 171586 136338 171822 136574
rect 171266 100658 171502 100894
rect 171586 100658 171822 100894
rect 171266 100338 171502 100574
rect 171586 100338 171822 100574
rect 171266 64658 171502 64894
rect 171586 64658 171822 64894
rect 171266 64338 171502 64574
rect 171586 64338 171822 64574
rect 171266 28658 171502 28894
rect 171586 28658 171822 28894
rect 171266 28338 171502 28574
rect 171586 28338 171822 28574
rect 171266 -5382 171502 -5146
rect 171586 -5382 171822 -5146
rect 171266 -5702 171502 -5466
rect 171586 -5702 171822 -5466
rect 174986 176378 175222 176614
rect 175306 176378 175542 176614
rect 174986 176058 175222 176294
rect 175306 176058 175542 176294
rect 174986 140378 175222 140614
rect 175306 140378 175542 140614
rect 174986 140058 175222 140294
rect 175306 140058 175542 140294
rect 174986 104378 175222 104614
rect 175306 104378 175542 104614
rect 174986 104058 175222 104294
rect 175306 104058 175542 104294
rect 174986 68378 175222 68614
rect 175306 68378 175542 68614
rect 174986 68058 175222 68294
rect 175306 68058 175542 68294
rect 174986 32378 175222 32614
rect 175306 32378 175542 32614
rect 174986 32058 175222 32294
rect 175306 32058 175542 32294
rect 156986 -6342 157222 -6106
rect 157306 -6342 157542 -6106
rect 156986 -6662 157222 -6426
rect 157306 -6662 157542 -6426
rect 181826 183218 182062 183454
rect 182146 183218 182382 183454
rect 181826 182898 182062 183134
rect 182146 182898 182382 183134
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 181826 111218 182062 111454
rect 182146 111218 182382 111454
rect 181826 110898 182062 111134
rect 182146 110898 182382 111134
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 185546 186938 185782 187174
rect 185866 186938 186102 187174
rect 185546 186618 185782 186854
rect 185866 186618 186102 186854
rect 185546 150938 185782 151174
rect 185866 150938 186102 151174
rect 185546 150618 185782 150854
rect 185866 150618 186102 150854
rect 185546 114938 185782 115174
rect 185866 114938 186102 115174
rect 185546 114618 185782 114854
rect 185866 114618 186102 114854
rect 185546 78938 185782 79174
rect 185866 78938 186102 79174
rect 185546 78618 185782 78854
rect 185866 78618 186102 78854
rect 185546 42938 185782 43174
rect 185866 42938 186102 43174
rect 185546 42618 185782 42854
rect 185866 42618 186102 42854
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 185546 -2502 185782 -2266
rect 185866 -2502 186102 -2266
rect 185546 -2822 185782 -2586
rect 185866 -2822 186102 -2586
rect 189266 190658 189502 190894
rect 189586 190658 189822 190894
rect 189266 190338 189502 190574
rect 189586 190338 189822 190574
rect 189266 154658 189502 154894
rect 189586 154658 189822 154894
rect 189266 154338 189502 154574
rect 189586 154338 189822 154574
rect 189266 118658 189502 118894
rect 189586 118658 189822 118894
rect 189266 118338 189502 118574
rect 189586 118338 189822 118574
rect 189266 82658 189502 82894
rect 189586 82658 189822 82894
rect 189266 82338 189502 82574
rect 189586 82338 189822 82574
rect 189266 46658 189502 46894
rect 189586 46658 189822 46894
rect 189266 46338 189502 46574
rect 189586 46338 189822 46574
rect 189266 10658 189502 10894
rect 189586 10658 189822 10894
rect 189266 10338 189502 10574
rect 189586 10338 189822 10574
rect 189266 -4422 189502 -4186
rect 189586 -4422 189822 -4186
rect 189266 -4742 189502 -4506
rect 189586 -4742 189822 -4506
rect 210986 711322 211222 711558
rect 211306 711322 211542 711558
rect 210986 711002 211222 711238
rect 211306 711002 211542 711238
rect 207266 709402 207502 709638
rect 207586 709402 207822 709638
rect 207266 709082 207502 709318
rect 207586 709082 207822 709318
rect 203546 707482 203782 707718
rect 203866 707482 204102 707718
rect 203546 707162 203782 707398
rect 203866 707162 204102 707398
rect 192986 698378 193222 698614
rect 193306 698378 193542 698614
rect 192986 698058 193222 698294
rect 193306 698058 193542 698294
rect 192986 662378 193222 662614
rect 193306 662378 193542 662614
rect 192986 662058 193222 662294
rect 193306 662058 193542 662294
rect 192986 626378 193222 626614
rect 193306 626378 193542 626614
rect 192986 626058 193222 626294
rect 193306 626058 193542 626294
rect 192986 590378 193222 590614
rect 193306 590378 193542 590614
rect 192986 590058 193222 590294
rect 193306 590058 193542 590294
rect 192986 554378 193222 554614
rect 193306 554378 193542 554614
rect 192986 554058 193222 554294
rect 193306 554058 193542 554294
rect 192986 518378 193222 518614
rect 193306 518378 193542 518614
rect 192986 518058 193222 518294
rect 193306 518058 193542 518294
rect 192986 482378 193222 482614
rect 193306 482378 193542 482614
rect 192986 482058 193222 482294
rect 193306 482058 193542 482294
rect 192986 446378 193222 446614
rect 193306 446378 193542 446614
rect 192986 446058 193222 446294
rect 193306 446058 193542 446294
rect 192986 410378 193222 410614
rect 193306 410378 193542 410614
rect 192986 410058 193222 410294
rect 193306 410058 193542 410294
rect 192986 374378 193222 374614
rect 193306 374378 193542 374614
rect 192986 374058 193222 374294
rect 193306 374058 193542 374294
rect 192986 338378 193222 338614
rect 193306 338378 193542 338614
rect 192986 338058 193222 338294
rect 193306 338058 193542 338294
rect 192986 302378 193222 302614
rect 193306 302378 193542 302614
rect 192986 302058 193222 302294
rect 193306 302058 193542 302294
rect 192986 266378 193222 266614
rect 193306 266378 193542 266614
rect 192986 266058 193222 266294
rect 193306 266058 193542 266294
rect 192986 230378 193222 230614
rect 193306 230378 193542 230614
rect 192986 230058 193222 230294
rect 193306 230058 193542 230294
rect 192986 194378 193222 194614
rect 193306 194378 193542 194614
rect 192986 194058 193222 194294
rect 193306 194058 193542 194294
rect 192986 158378 193222 158614
rect 193306 158378 193542 158614
rect 192986 158058 193222 158294
rect 193306 158058 193542 158294
rect 192986 122378 193222 122614
rect 193306 122378 193542 122614
rect 192986 122058 193222 122294
rect 193306 122058 193542 122294
rect 192986 86378 193222 86614
rect 193306 86378 193542 86614
rect 192986 86058 193222 86294
rect 193306 86058 193542 86294
rect 192986 50378 193222 50614
rect 193306 50378 193542 50614
rect 192986 50058 193222 50294
rect 193306 50058 193542 50294
rect 192986 14378 193222 14614
rect 193306 14378 193542 14614
rect 192986 14058 193222 14294
rect 193306 14058 193542 14294
rect 174986 -7302 175222 -7066
rect 175306 -7302 175542 -7066
rect 174986 -7622 175222 -7386
rect 175306 -7622 175542 -7386
rect 199826 705562 200062 705798
rect 200146 705562 200382 705798
rect 199826 705242 200062 705478
rect 200146 705242 200382 705478
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 199826 561218 200062 561454
rect 200146 561218 200382 561454
rect 199826 560898 200062 561134
rect 200146 560898 200382 561134
rect 199826 525218 200062 525454
rect 200146 525218 200382 525454
rect 199826 524898 200062 525134
rect 200146 524898 200382 525134
rect 199826 489218 200062 489454
rect 200146 489218 200382 489454
rect 199826 488898 200062 489134
rect 200146 488898 200382 489134
rect 199826 453218 200062 453454
rect 200146 453218 200382 453454
rect 199826 452898 200062 453134
rect 200146 452898 200382 453134
rect 199826 417218 200062 417454
rect 200146 417218 200382 417454
rect 199826 416898 200062 417134
rect 200146 416898 200382 417134
rect 199826 381218 200062 381454
rect 200146 381218 200382 381454
rect 199826 380898 200062 381134
rect 200146 380898 200382 381134
rect 199826 345218 200062 345454
rect 200146 345218 200382 345454
rect 199826 344898 200062 345134
rect 200146 344898 200382 345134
rect 199826 309218 200062 309454
rect 200146 309218 200382 309454
rect 199826 308898 200062 309134
rect 200146 308898 200382 309134
rect 199826 273218 200062 273454
rect 200146 273218 200382 273454
rect 199826 272898 200062 273134
rect 200146 272898 200382 273134
rect 199826 237218 200062 237454
rect 200146 237218 200382 237454
rect 199826 236898 200062 237134
rect 200146 236898 200382 237134
rect 199826 201218 200062 201454
rect 200146 201218 200382 201454
rect 199826 200898 200062 201134
rect 200146 200898 200382 201134
rect 199826 165218 200062 165454
rect 200146 165218 200382 165454
rect 199826 164898 200062 165134
rect 200146 164898 200382 165134
rect 199826 129218 200062 129454
rect 200146 129218 200382 129454
rect 199826 128898 200062 129134
rect 200146 128898 200382 129134
rect 199826 93218 200062 93454
rect 200146 93218 200382 93454
rect 199826 92898 200062 93134
rect 200146 92898 200382 93134
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -1542 200062 -1306
rect 200146 -1542 200382 -1306
rect 199826 -1862 200062 -1626
rect 200146 -1862 200382 -1626
rect 203546 672938 203782 673174
rect 203866 672938 204102 673174
rect 203546 672618 203782 672854
rect 203866 672618 204102 672854
rect 203546 636938 203782 637174
rect 203866 636938 204102 637174
rect 203546 636618 203782 636854
rect 203866 636618 204102 636854
rect 203546 600938 203782 601174
rect 203866 600938 204102 601174
rect 203546 600618 203782 600854
rect 203866 600618 204102 600854
rect 203546 564938 203782 565174
rect 203866 564938 204102 565174
rect 203546 564618 203782 564854
rect 203866 564618 204102 564854
rect 203546 528938 203782 529174
rect 203866 528938 204102 529174
rect 203546 528618 203782 528854
rect 203866 528618 204102 528854
rect 203546 492938 203782 493174
rect 203866 492938 204102 493174
rect 203546 492618 203782 492854
rect 203866 492618 204102 492854
rect 203546 456938 203782 457174
rect 203866 456938 204102 457174
rect 203546 456618 203782 456854
rect 203866 456618 204102 456854
rect 203546 420938 203782 421174
rect 203866 420938 204102 421174
rect 203546 420618 203782 420854
rect 203866 420618 204102 420854
rect 203546 384938 203782 385174
rect 203866 384938 204102 385174
rect 203546 384618 203782 384854
rect 203866 384618 204102 384854
rect 203546 348938 203782 349174
rect 203866 348938 204102 349174
rect 203546 348618 203782 348854
rect 203866 348618 204102 348854
rect 203546 312938 203782 313174
rect 203866 312938 204102 313174
rect 203546 312618 203782 312854
rect 203866 312618 204102 312854
rect 203546 276938 203782 277174
rect 203866 276938 204102 277174
rect 203546 276618 203782 276854
rect 203866 276618 204102 276854
rect 203546 240938 203782 241174
rect 203866 240938 204102 241174
rect 203546 240618 203782 240854
rect 203866 240618 204102 240854
rect 203546 204938 203782 205174
rect 203866 204938 204102 205174
rect 203546 204618 203782 204854
rect 203866 204618 204102 204854
rect 203546 168938 203782 169174
rect 203866 168938 204102 169174
rect 203546 168618 203782 168854
rect 203866 168618 204102 168854
rect 203546 132938 203782 133174
rect 203866 132938 204102 133174
rect 203546 132618 203782 132854
rect 203866 132618 204102 132854
rect 203546 96938 203782 97174
rect 203866 96938 204102 97174
rect 203546 96618 203782 96854
rect 203866 96618 204102 96854
rect 203546 60938 203782 61174
rect 203866 60938 204102 61174
rect 203546 60618 203782 60854
rect 203866 60618 204102 60854
rect 203546 24938 203782 25174
rect 203866 24938 204102 25174
rect 203546 24618 203782 24854
rect 203866 24618 204102 24854
rect 203546 -3462 203782 -3226
rect 203866 -3462 204102 -3226
rect 203546 -3782 203782 -3546
rect 203866 -3782 204102 -3546
rect 207266 676658 207502 676894
rect 207586 676658 207822 676894
rect 207266 676338 207502 676574
rect 207586 676338 207822 676574
rect 207266 640658 207502 640894
rect 207586 640658 207822 640894
rect 207266 640338 207502 640574
rect 207586 640338 207822 640574
rect 207266 604658 207502 604894
rect 207586 604658 207822 604894
rect 207266 604338 207502 604574
rect 207586 604338 207822 604574
rect 207266 568658 207502 568894
rect 207586 568658 207822 568894
rect 207266 568338 207502 568574
rect 207586 568338 207822 568574
rect 207266 532658 207502 532894
rect 207586 532658 207822 532894
rect 207266 532338 207502 532574
rect 207586 532338 207822 532574
rect 207266 496658 207502 496894
rect 207586 496658 207822 496894
rect 207266 496338 207502 496574
rect 207586 496338 207822 496574
rect 207266 460658 207502 460894
rect 207586 460658 207822 460894
rect 207266 460338 207502 460574
rect 207586 460338 207822 460574
rect 207266 424658 207502 424894
rect 207586 424658 207822 424894
rect 207266 424338 207502 424574
rect 207586 424338 207822 424574
rect 207266 388658 207502 388894
rect 207586 388658 207822 388894
rect 207266 388338 207502 388574
rect 207586 388338 207822 388574
rect 207266 352658 207502 352894
rect 207586 352658 207822 352894
rect 207266 352338 207502 352574
rect 207586 352338 207822 352574
rect 207266 316658 207502 316894
rect 207586 316658 207822 316894
rect 207266 316338 207502 316574
rect 207586 316338 207822 316574
rect 207266 280658 207502 280894
rect 207586 280658 207822 280894
rect 207266 280338 207502 280574
rect 207586 280338 207822 280574
rect 207266 244658 207502 244894
rect 207586 244658 207822 244894
rect 207266 244338 207502 244574
rect 207586 244338 207822 244574
rect 207266 208658 207502 208894
rect 207586 208658 207822 208894
rect 207266 208338 207502 208574
rect 207586 208338 207822 208574
rect 207266 172658 207502 172894
rect 207586 172658 207822 172894
rect 207266 172338 207502 172574
rect 207586 172338 207822 172574
rect 207266 136658 207502 136894
rect 207586 136658 207822 136894
rect 207266 136338 207502 136574
rect 207586 136338 207822 136574
rect 207266 100658 207502 100894
rect 207586 100658 207822 100894
rect 207266 100338 207502 100574
rect 207586 100338 207822 100574
rect 207266 64658 207502 64894
rect 207586 64658 207822 64894
rect 207266 64338 207502 64574
rect 207586 64338 207822 64574
rect 207266 28658 207502 28894
rect 207586 28658 207822 28894
rect 207266 28338 207502 28574
rect 207586 28338 207822 28574
rect 207266 -5382 207502 -5146
rect 207586 -5382 207822 -5146
rect 207266 -5702 207502 -5466
rect 207586 -5702 207822 -5466
rect 228986 710362 229222 710598
rect 229306 710362 229542 710598
rect 228986 710042 229222 710278
rect 229306 710042 229542 710278
rect 225266 708442 225502 708678
rect 225586 708442 225822 708678
rect 225266 708122 225502 708358
rect 225586 708122 225822 708358
rect 221546 706522 221782 706758
rect 221866 706522 222102 706758
rect 221546 706202 221782 706438
rect 221866 706202 222102 706438
rect 210986 680378 211222 680614
rect 211306 680378 211542 680614
rect 210986 680058 211222 680294
rect 211306 680058 211542 680294
rect 210986 644378 211222 644614
rect 211306 644378 211542 644614
rect 210986 644058 211222 644294
rect 211306 644058 211542 644294
rect 210986 608378 211222 608614
rect 211306 608378 211542 608614
rect 210986 608058 211222 608294
rect 211306 608058 211542 608294
rect 210986 572378 211222 572614
rect 211306 572378 211542 572614
rect 210986 572058 211222 572294
rect 211306 572058 211542 572294
rect 210986 536378 211222 536614
rect 211306 536378 211542 536614
rect 210986 536058 211222 536294
rect 211306 536058 211542 536294
rect 210986 500378 211222 500614
rect 211306 500378 211542 500614
rect 210986 500058 211222 500294
rect 211306 500058 211542 500294
rect 210986 464378 211222 464614
rect 211306 464378 211542 464614
rect 210986 464058 211222 464294
rect 211306 464058 211542 464294
rect 210986 428378 211222 428614
rect 211306 428378 211542 428614
rect 210986 428058 211222 428294
rect 211306 428058 211542 428294
rect 210986 392378 211222 392614
rect 211306 392378 211542 392614
rect 210986 392058 211222 392294
rect 211306 392058 211542 392294
rect 210986 356378 211222 356614
rect 211306 356378 211542 356614
rect 210986 356058 211222 356294
rect 211306 356058 211542 356294
rect 210986 320378 211222 320614
rect 211306 320378 211542 320614
rect 210986 320058 211222 320294
rect 211306 320058 211542 320294
rect 210986 284378 211222 284614
rect 211306 284378 211542 284614
rect 210986 284058 211222 284294
rect 211306 284058 211542 284294
rect 210986 248378 211222 248614
rect 211306 248378 211542 248614
rect 210986 248058 211222 248294
rect 211306 248058 211542 248294
rect 210986 212378 211222 212614
rect 211306 212378 211542 212614
rect 210986 212058 211222 212294
rect 211306 212058 211542 212294
rect 210986 176378 211222 176614
rect 211306 176378 211542 176614
rect 210986 176058 211222 176294
rect 211306 176058 211542 176294
rect 210986 140378 211222 140614
rect 211306 140378 211542 140614
rect 210986 140058 211222 140294
rect 211306 140058 211542 140294
rect 210986 104378 211222 104614
rect 211306 104378 211542 104614
rect 210986 104058 211222 104294
rect 211306 104058 211542 104294
rect 210986 68378 211222 68614
rect 211306 68378 211542 68614
rect 210986 68058 211222 68294
rect 211306 68058 211542 68294
rect 210986 32378 211222 32614
rect 211306 32378 211542 32614
rect 210986 32058 211222 32294
rect 211306 32058 211542 32294
rect 192986 -6342 193222 -6106
rect 193306 -6342 193542 -6106
rect 192986 -6662 193222 -6426
rect 193306 -6662 193542 -6426
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 217826 543218 218062 543454
rect 218146 543218 218382 543454
rect 217826 542898 218062 543134
rect 218146 542898 218382 543134
rect 217826 507218 218062 507454
rect 218146 507218 218382 507454
rect 217826 506898 218062 507134
rect 218146 506898 218382 507134
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 217826 435218 218062 435454
rect 218146 435218 218382 435454
rect 217826 434898 218062 435134
rect 218146 434898 218382 435134
rect 217826 399218 218062 399454
rect 218146 399218 218382 399454
rect 217826 398898 218062 399134
rect 218146 398898 218382 399134
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 217826 327218 218062 327454
rect 218146 327218 218382 327454
rect 217826 326898 218062 327134
rect 218146 326898 218382 327134
rect 217826 291218 218062 291454
rect 218146 291218 218382 291454
rect 217826 290898 218062 291134
rect 218146 290898 218382 291134
rect 217826 255218 218062 255454
rect 218146 255218 218382 255454
rect 217826 254898 218062 255134
rect 218146 254898 218382 255134
rect 217826 219218 218062 219454
rect 218146 219218 218382 219454
rect 217826 218898 218062 219134
rect 218146 218898 218382 219134
rect 217826 183218 218062 183454
rect 218146 183218 218382 183454
rect 217826 182898 218062 183134
rect 218146 182898 218382 183134
rect 217826 147218 218062 147454
rect 218146 147218 218382 147454
rect 217826 146898 218062 147134
rect 218146 146898 218382 147134
rect 217826 111218 218062 111454
rect 218146 111218 218382 111454
rect 217826 110898 218062 111134
rect 218146 110898 218382 111134
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 221546 690938 221782 691174
rect 221866 690938 222102 691174
rect 221546 690618 221782 690854
rect 221866 690618 222102 690854
rect 221546 654938 221782 655174
rect 221866 654938 222102 655174
rect 221546 654618 221782 654854
rect 221866 654618 222102 654854
rect 221546 618938 221782 619174
rect 221866 618938 222102 619174
rect 221546 618618 221782 618854
rect 221866 618618 222102 618854
rect 221546 582938 221782 583174
rect 221866 582938 222102 583174
rect 221546 582618 221782 582854
rect 221866 582618 222102 582854
rect 221546 546938 221782 547174
rect 221866 546938 222102 547174
rect 221546 546618 221782 546854
rect 221866 546618 222102 546854
rect 221546 510938 221782 511174
rect 221866 510938 222102 511174
rect 221546 510618 221782 510854
rect 221866 510618 222102 510854
rect 221546 474938 221782 475174
rect 221866 474938 222102 475174
rect 221546 474618 221782 474854
rect 221866 474618 222102 474854
rect 221546 438938 221782 439174
rect 221866 438938 222102 439174
rect 221546 438618 221782 438854
rect 221866 438618 222102 438854
rect 221546 402938 221782 403174
rect 221866 402938 222102 403174
rect 221546 402618 221782 402854
rect 221866 402618 222102 402854
rect 221546 366938 221782 367174
rect 221866 366938 222102 367174
rect 221546 366618 221782 366854
rect 221866 366618 222102 366854
rect 221546 330938 221782 331174
rect 221866 330938 222102 331174
rect 221546 330618 221782 330854
rect 221866 330618 222102 330854
rect 221546 294938 221782 295174
rect 221866 294938 222102 295174
rect 221546 294618 221782 294854
rect 221866 294618 222102 294854
rect 221546 258938 221782 259174
rect 221866 258938 222102 259174
rect 221546 258618 221782 258854
rect 221866 258618 222102 258854
rect 221546 222938 221782 223174
rect 221866 222938 222102 223174
rect 221546 222618 221782 222854
rect 221866 222618 222102 222854
rect 221546 186938 221782 187174
rect 221866 186938 222102 187174
rect 221546 186618 221782 186854
rect 221866 186618 222102 186854
rect 221546 150938 221782 151174
rect 221866 150938 222102 151174
rect 221546 150618 221782 150854
rect 221866 150618 222102 150854
rect 221546 114938 221782 115174
rect 221866 114938 222102 115174
rect 221546 114618 221782 114854
rect 221866 114618 222102 114854
rect 221546 78938 221782 79174
rect 221866 78938 222102 79174
rect 221546 78618 221782 78854
rect 221866 78618 222102 78854
rect 221546 42938 221782 43174
rect 221866 42938 222102 43174
rect 221546 42618 221782 42854
rect 221866 42618 222102 42854
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 221546 -2502 221782 -2266
rect 221866 -2502 222102 -2266
rect 221546 -2822 221782 -2586
rect 221866 -2822 222102 -2586
rect 225266 694658 225502 694894
rect 225586 694658 225822 694894
rect 225266 694338 225502 694574
rect 225586 694338 225822 694574
rect 225266 658658 225502 658894
rect 225586 658658 225822 658894
rect 225266 658338 225502 658574
rect 225586 658338 225822 658574
rect 225266 622658 225502 622894
rect 225586 622658 225822 622894
rect 225266 622338 225502 622574
rect 225586 622338 225822 622574
rect 225266 586658 225502 586894
rect 225586 586658 225822 586894
rect 225266 586338 225502 586574
rect 225586 586338 225822 586574
rect 225266 550658 225502 550894
rect 225586 550658 225822 550894
rect 225266 550338 225502 550574
rect 225586 550338 225822 550574
rect 225266 514658 225502 514894
rect 225586 514658 225822 514894
rect 225266 514338 225502 514574
rect 225586 514338 225822 514574
rect 225266 478658 225502 478894
rect 225586 478658 225822 478894
rect 225266 478338 225502 478574
rect 225586 478338 225822 478574
rect 225266 442658 225502 442894
rect 225586 442658 225822 442894
rect 225266 442338 225502 442574
rect 225586 442338 225822 442574
rect 225266 406658 225502 406894
rect 225586 406658 225822 406894
rect 225266 406338 225502 406574
rect 225586 406338 225822 406574
rect 225266 370658 225502 370894
rect 225586 370658 225822 370894
rect 225266 370338 225502 370574
rect 225586 370338 225822 370574
rect 225266 334658 225502 334894
rect 225586 334658 225822 334894
rect 225266 334338 225502 334574
rect 225586 334338 225822 334574
rect 225266 298658 225502 298894
rect 225586 298658 225822 298894
rect 225266 298338 225502 298574
rect 225586 298338 225822 298574
rect 225266 262658 225502 262894
rect 225586 262658 225822 262894
rect 225266 262338 225502 262574
rect 225586 262338 225822 262574
rect 225266 226658 225502 226894
rect 225586 226658 225822 226894
rect 225266 226338 225502 226574
rect 225586 226338 225822 226574
rect 225266 190658 225502 190894
rect 225586 190658 225822 190894
rect 225266 190338 225502 190574
rect 225586 190338 225822 190574
rect 225266 154658 225502 154894
rect 225586 154658 225822 154894
rect 225266 154338 225502 154574
rect 225586 154338 225822 154574
rect 225266 118658 225502 118894
rect 225586 118658 225822 118894
rect 225266 118338 225502 118574
rect 225586 118338 225822 118574
rect 225266 82658 225502 82894
rect 225586 82658 225822 82894
rect 225266 82338 225502 82574
rect 225586 82338 225822 82574
rect 225266 46658 225502 46894
rect 225586 46658 225822 46894
rect 225266 46338 225502 46574
rect 225586 46338 225822 46574
rect 225266 10658 225502 10894
rect 225586 10658 225822 10894
rect 225266 10338 225502 10574
rect 225586 10338 225822 10574
rect 225266 -4422 225502 -4186
rect 225586 -4422 225822 -4186
rect 225266 -4742 225502 -4506
rect 225586 -4742 225822 -4506
rect 246986 711322 247222 711558
rect 247306 711322 247542 711558
rect 246986 711002 247222 711238
rect 247306 711002 247542 711238
rect 243266 709402 243502 709638
rect 243586 709402 243822 709638
rect 243266 709082 243502 709318
rect 243586 709082 243822 709318
rect 239546 707482 239782 707718
rect 239866 707482 240102 707718
rect 239546 707162 239782 707398
rect 239866 707162 240102 707398
rect 235826 705562 236062 705798
rect 236146 705562 236382 705798
rect 235826 705242 236062 705478
rect 236146 705242 236382 705478
rect 228986 698378 229222 698614
rect 229306 698378 229542 698614
rect 228986 698058 229222 698294
rect 229306 698058 229542 698294
rect 228986 662378 229222 662614
rect 229306 662378 229542 662614
rect 228986 662058 229222 662294
rect 229306 662058 229542 662294
rect 228986 626378 229222 626614
rect 229306 626378 229542 626614
rect 228986 626058 229222 626294
rect 229306 626058 229542 626294
rect 228986 590378 229222 590614
rect 229306 590378 229542 590614
rect 228986 590058 229222 590294
rect 229306 590058 229542 590294
rect 228986 554378 229222 554614
rect 229306 554378 229542 554614
rect 228986 554058 229222 554294
rect 229306 554058 229542 554294
rect 228986 518378 229222 518614
rect 229306 518378 229542 518614
rect 228986 518058 229222 518294
rect 229306 518058 229542 518294
rect 228986 482378 229222 482614
rect 229306 482378 229542 482614
rect 228986 482058 229222 482294
rect 229306 482058 229542 482294
rect 228986 446378 229222 446614
rect 229306 446378 229542 446614
rect 228986 446058 229222 446294
rect 229306 446058 229542 446294
rect 228986 410378 229222 410614
rect 229306 410378 229542 410614
rect 228986 410058 229222 410294
rect 229306 410058 229542 410294
rect 228986 374378 229222 374614
rect 229306 374378 229542 374614
rect 228986 374058 229222 374294
rect 229306 374058 229542 374294
rect 228986 338378 229222 338614
rect 229306 338378 229542 338614
rect 228986 338058 229222 338294
rect 229306 338058 229542 338294
rect 228986 302378 229222 302614
rect 229306 302378 229542 302614
rect 228986 302058 229222 302294
rect 229306 302058 229542 302294
rect 228986 266378 229222 266614
rect 229306 266378 229542 266614
rect 228986 266058 229222 266294
rect 229306 266058 229542 266294
rect 228986 230378 229222 230614
rect 229306 230378 229542 230614
rect 228986 230058 229222 230294
rect 229306 230058 229542 230294
rect 228986 194378 229222 194614
rect 229306 194378 229542 194614
rect 228986 194058 229222 194294
rect 229306 194058 229542 194294
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 235826 561218 236062 561454
rect 236146 561218 236382 561454
rect 235826 560898 236062 561134
rect 236146 560898 236382 561134
rect 235826 525218 236062 525454
rect 236146 525218 236382 525454
rect 235826 524898 236062 525134
rect 236146 524898 236382 525134
rect 235826 489218 236062 489454
rect 236146 489218 236382 489454
rect 235826 488898 236062 489134
rect 236146 488898 236382 489134
rect 235826 453218 236062 453454
rect 236146 453218 236382 453454
rect 235826 452898 236062 453134
rect 236146 452898 236382 453134
rect 235826 417218 236062 417454
rect 236146 417218 236382 417454
rect 235826 416898 236062 417134
rect 236146 416898 236382 417134
rect 235826 381218 236062 381454
rect 236146 381218 236382 381454
rect 235826 380898 236062 381134
rect 236146 380898 236382 381134
rect 235826 345218 236062 345454
rect 236146 345218 236382 345454
rect 235826 344898 236062 345134
rect 236146 344898 236382 345134
rect 235826 309218 236062 309454
rect 236146 309218 236382 309454
rect 235826 308898 236062 309134
rect 236146 308898 236382 309134
rect 235826 273218 236062 273454
rect 236146 273218 236382 273454
rect 235826 272898 236062 273134
rect 236146 272898 236382 273134
rect 235826 237218 236062 237454
rect 236146 237218 236382 237454
rect 235826 236898 236062 237134
rect 236146 236898 236382 237134
rect 235826 201218 236062 201454
rect 236146 201218 236382 201454
rect 235826 200898 236062 201134
rect 236146 200898 236382 201134
rect 228986 158378 229222 158614
rect 229306 158378 229542 158614
rect 228986 158058 229222 158294
rect 229306 158058 229542 158294
rect 228986 122378 229222 122614
rect 229306 122378 229542 122614
rect 228986 122058 229222 122294
rect 229306 122058 229542 122294
rect 228986 86378 229222 86614
rect 229306 86378 229542 86614
rect 228986 86058 229222 86294
rect 229306 86058 229542 86294
rect 228986 50378 229222 50614
rect 229306 50378 229542 50614
rect 228986 50058 229222 50294
rect 229306 50058 229542 50294
rect 228986 14378 229222 14614
rect 229306 14378 229542 14614
rect 228986 14058 229222 14294
rect 229306 14058 229542 14294
rect 210986 -7302 211222 -7066
rect 211306 -7302 211542 -7066
rect 210986 -7622 211222 -7386
rect 211306 -7622 211542 -7386
rect 239546 672938 239782 673174
rect 239866 672938 240102 673174
rect 239546 672618 239782 672854
rect 239866 672618 240102 672854
rect 239546 636938 239782 637174
rect 239866 636938 240102 637174
rect 239546 636618 239782 636854
rect 239866 636618 240102 636854
rect 239546 600938 239782 601174
rect 239866 600938 240102 601174
rect 239546 600618 239782 600854
rect 239866 600618 240102 600854
rect 239546 564938 239782 565174
rect 239866 564938 240102 565174
rect 239546 564618 239782 564854
rect 239866 564618 240102 564854
rect 239546 528938 239782 529174
rect 239866 528938 240102 529174
rect 239546 528618 239782 528854
rect 239866 528618 240102 528854
rect 239546 492938 239782 493174
rect 239866 492938 240102 493174
rect 239546 492618 239782 492854
rect 239866 492618 240102 492854
rect 243266 676658 243502 676894
rect 243586 676658 243822 676894
rect 243266 676338 243502 676574
rect 243586 676338 243822 676574
rect 243266 640658 243502 640894
rect 243586 640658 243822 640894
rect 243266 640338 243502 640574
rect 243586 640338 243822 640574
rect 243266 604658 243502 604894
rect 243586 604658 243822 604894
rect 243266 604338 243502 604574
rect 243586 604338 243822 604574
rect 243266 568658 243502 568894
rect 243586 568658 243822 568894
rect 243266 568338 243502 568574
rect 243586 568338 243822 568574
rect 243266 532658 243502 532894
rect 243586 532658 243822 532894
rect 243266 532338 243502 532574
rect 243586 532338 243822 532574
rect 243266 496658 243502 496894
rect 243586 496658 243822 496894
rect 243266 496338 243502 496574
rect 243586 496338 243822 496574
rect 264986 710362 265222 710598
rect 265306 710362 265542 710598
rect 264986 710042 265222 710278
rect 265306 710042 265542 710278
rect 261266 708442 261502 708678
rect 261586 708442 261822 708678
rect 261266 708122 261502 708358
rect 261586 708122 261822 708358
rect 257546 706522 257782 706758
rect 257866 706522 258102 706758
rect 257546 706202 257782 706438
rect 257866 706202 258102 706438
rect 246986 680378 247222 680614
rect 247306 680378 247542 680614
rect 246986 680058 247222 680294
rect 247306 680058 247542 680294
rect 246986 644378 247222 644614
rect 247306 644378 247542 644614
rect 246986 644058 247222 644294
rect 247306 644058 247542 644294
rect 246986 608378 247222 608614
rect 247306 608378 247542 608614
rect 246986 608058 247222 608294
rect 247306 608058 247542 608294
rect 246986 572378 247222 572614
rect 247306 572378 247542 572614
rect 246986 572058 247222 572294
rect 247306 572058 247542 572294
rect 246986 536378 247222 536614
rect 247306 536378 247542 536614
rect 246986 536058 247222 536294
rect 247306 536058 247542 536294
rect 246986 500378 247222 500614
rect 247306 500378 247542 500614
rect 246986 500058 247222 500294
rect 247306 500058 247542 500294
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 253826 543218 254062 543454
rect 254146 543218 254382 543454
rect 253826 542898 254062 543134
rect 254146 542898 254382 543134
rect 253826 507218 254062 507454
rect 254146 507218 254382 507454
rect 253826 506898 254062 507134
rect 254146 506898 254382 507134
rect 257546 690938 257782 691174
rect 257866 690938 258102 691174
rect 257546 690618 257782 690854
rect 257866 690618 258102 690854
rect 257546 654938 257782 655174
rect 257866 654938 258102 655174
rect 257546 654618 257782 654854
rect 257866 654618 258102 654854
rect 257546 618938 257782 619174
rect 257866 618938 258102 619174
rect 257546 618618 257782 618854
rect 257866 618618 258102 618854
rect 257546 582938 257782 583174
rect 257866 582938 258102 583174
rect 257546 582618 257782 582854
rect 257866 582618 258102 582854
rect 257546 546938 257782 547174
rect 257866 546938 258102 547174
rect 257546 546618 257782 546854
rect 257866 546618 258102 546854
rect 257546 510938 257782 511174
rect 257866 510938 258102 511174
rect 257546 510618 257782 510854
rect 257866 510618 258102 510854
rect 261266 694658 261502 694894
rect 261586 694658 261822 694894
rect 261266 694338 261502 694574
rect 261586 694338 261822 694574
rect 261266 658658 261502 658894
rect 261586 658658 261822 658894
rect 261266 658338 261502 658574
rect 261586 658338 261822 658574
rect 261266 622658 261502 622894
rect 261586 622658 261822 622894
rect 261266 622338 261502 622574
rect 261586 622338 261822 622574
rect 261266 586658 261502 586894
rect 261586 586658 261822 586894
rect 261266 586338 261502 586574
rect 261586 586338 261822 586574
rect 261266 550658 261502 550894
rect 261586 550658 261822 550894
rect 261266 550338 261502 550574
rect 261586 550338 261822 550574
rect 261266 514658 261502 514894
rect 261586 514658 261822 514894
rect 261266 514338 261502 514574
rect 261586 514338 261822 514574
rect 282986 711322 283222 711558
rect 283306 711322 283542 711558
rect 282986 711002 283222 711238
rect 283306 711002 283542 711238
rect 279266 709402 279502 709638
rect 279586 709402 279822 709638
rect 279266 709082 279502 709318
rect 279586 709082 279822 709318
rect 275546 707482 275782 707718
rect 275866 707482 276102 707718
rect 275546 707162 275782 707398
rect 275866 707162 276102 707398
rect 264986 698378 265222 698614
rect 265306 698378 265542 698614
rect 264986 698058 265222 698294
rect 265306 698058 265542 698294
rect 264986 662378 265222 662614
rect 265306 662378 265542 662614
rect 264986 662058 265222 662294
rect 265306 662058 265542 662294
rect 264986 626378 265222 626614
rect 265306 626378 265542 626614
rect 264986 626058 265222 626294
rect 265306 626058 265542 626294
rect 264986 590378 265222 590614
rect 265306 590378 265542 590614
rect 264986 590058 265222 590294
rect 265306 590058 265542 590294
rect 264986 554378 265222 554614
rect 265306 554378 265542 554614
rect 264986 554058 265222 554294
rect 265306 554058 265542 554294
rect 264986 518378 265222 518614
rect 265306 518378 265542 518614
rect 264986 518058 265222 518294
rect 265306 518058 265542 518294
rect 264986 482378 265222 482614
rect 265306 482378 265542 482614
rect 264986 482058 265222 482294
rect 265306 482058 265542 482294
rect 271826 705562 272062 705798
rect 272146 705562 272382 705798
rect 271826 705242 272062 705478
rect 272146 705242 272382 705478
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 271826 561218 272062 561454
rect 272146 561218 272382 561454
rect 271826 560898 272062 561134
rect 272146 560898 272382 561134
rect 271826 525218 272062 525454
rect 272146 525218 272382 525454
rect 271826 524898 272062 525134
rect 272146 524898 272382 525134
rect 271826 489218 272062 489454
rect 272146 489218 272382 489454
rect 271826 488898 272062 489134
rect 272146 488898 272382 489134
rect 275546 672938 275782 673174
rect 275866 672938 276102 673174
rect 275546 672618 275782 672854
rect 275866 672618 276102 672854
rect 275546 636938 275782 637174
rect 275866 636938 276102 637174
rect 275546 636618 275782 636854
rect 275866 636618 276102 636854
rect 275546 600938 275782 601174
rect 275866 600938 276102 601174
rect 275546 600618 275782 600854
rect 275866 600618 276102 600854
rect 275546 564938 275782 565174
rect 275866 564938 276102 565174
rect 275546 564618 275782 564854
rect 275866 564618 276102 564854
rect 275546 528938 275782 529174
rect 275866 528938 276102 529174
rect 275546 528618 275782 528854
rect 275866 528618 276102 528854
rect 275546 492938 275782 493174
rect 275866 492938 276102 493174
rect 275546 492618 275782 492854
rect 275866 492618 276102 492854
rect 279266 676658 279502 676894
rect 279586 676658 279822 676894
rect 279266 676338 279502 676574
rect 279586 676338 279822 676574
rect 279266 640658 279502 640894
rect 279586 640658 279822 640894
rect 279266 640338 279502 640574
rect 279586 640338 279822 640574
rect 279266 604658 279502 604894
rect 279586 604658 279822 604894
rect 279266 604338 279502 604574
rect 279586 604338 279822 604574
rect 279266 568658 279502 568894
rect 279586 568658 279822 568894
rect 279266 568338 279502 568574
rect 279586 568338 279822 568574
rect 279266 532658 279502 532894
rect 279586 532658 279822 532894
rect 279266 532338 279502 532574
rect 279586 532338 279822 532574
rect 279266 496658 279502 496894
rect 279586 496658 279822 496894
rect 279266 496338 279502 496574
rect 279586 496338 279822 496574
rect 300986 710362 301222 710598
rect 301306 710362 301542 710598
rect 300986 710042 301222 710278
rect 301306 710042 301542 710278
rect 297266 708442 297502 708678
rect 297586 708442 297822 708678
rect 297266 708122 297502 708358
rect 297586 708122 297822 708358
rect 293546 706522 293782 706758
rect 293866 706522 294102 706758
rect 293546 706202 293782 706438
rect 293866 706202 294102 706438
rect 282986 680378 283222 680614
rect 283306 680378 283542 680614
rect 282986 680058 283222 680294
rect 283306 680058 283542 680294
rect 282986 644378 283222 644614
rect 283306 644378 283542 644614
rect 282986 644058 283222 644294
rect 283306 644058 283542 644294
rect 282986 608378 283222 608614
rect 283306 608378 283542 608614
rect 282986 608058 283222 608294
rect 283306 608058 283542 608294
rect 282986 572378 283222 572614
rect 283306 572378 283542 572614
rect 282986 572058 283222 572294
rect 283306 572058 283542 572294
rect 282986 536378 283222 536614
rect 283306 536378 283542 536614
rect 282986 536058 283222 536294
rect 283306 536058 283542 536294
rect 282986 500378 283222 500614
rect 283306 500378 283542 500614
rect 282986 500058 283222 500294
rect 283306 500058 283542 500294
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 289826 507218 290062 507454
rect 290146 507218 290382 507454
rect 289826 506898 290062 507134
rect 290146 506898 290382 507134
rect 293546 690938 293782 691174
rect 293866 690938 294102 691174
rect 293546 690618 293782 690854
rect 293866 690618 294102 690854
rect 293546 654938 293782 655174
rect 293866 654938 294102 655174
rect 293546 654618 293782 654854
rect 293866 654618 294102 654854
rect 293546 618938 293782 619174
rect 293866 618938 294102 619174
rect 293546 618618 293782 618854
rect 293866 618618 294102 618854
rect 293546 582938 293782 583174
rect 293866 582938 294102 583174
rect 293546 582618 293782 582854
rect 293866 582618 294102 582854
rect 293546 546938 293782 547174
rect 293866 546938 294102 547174
rect 293546 546618 293782 546854
rect 293866 546618 294102 546854
rect 293546 510938 293782 511174
rect 293866 510938 294102 511174
rect 293546 510618 293782 510854
rect 293866 510618 294102 510854
rect 297266 694658 297502 694894
rect 297586 694658 297822 694894
rect 297266 694338 297502 694574
rect 297586 694338 297822 694574
rect 297266 658658 297502 658894
rect 297586 658658 297822 658894
rect 297266 658338 297502 658574
rect 297586 658338 297822 658574
rect 297266 622658 297502 622894
rect 297586 622658 297822 622894
rect 297266 622338 297502 622574
rect 297586 622338 297822 622574
rect 297266 586658 297502 586894
rect 297586 586658 297822 586894
rect 297266 586338 297502 586574
rect 297586 586338 297822 586574
rect 297266 550658 297502 550894
rect 297586 550658 297822 550894
rect 297266 550338 297502 550574
rect 297586 550338 297822 550574
rect 297266 514658 297502 514894
rect 297586 514658 297822 514894
rect 297266 514338 297502 514574
rect 297586 514338 297822 514574
rect 318986 711322 319222 711558
rect 319306 711322 319542 711558
rect 318986 711002 319222 711238
rect 319306 711002 319542 711238
rect 315266 709402 315502 709638
rect 315586 709402 315822 709638
rect 315266 709082 315502 709318
rect 315586 709082 315822 709318
rect 311546 707482 311782 707718
rect 311866 707482 312102 707718
rect 311546 707162 311782 707398
rect 311866 707162 312102 707398
rect 300986 698378 301222 698614
rect 301306 698378 301542 698614
rect 300986 698058 301222 698294
rect 301306 698058 301542 698294
rect 300986 662378 301222 662614
rect 301306 662378 301542 662614
rect 300986 662058 301222 662294
rect 301306 662058 301542 662294
rect 300986 626378 301222 626614
rect 301306 626378 301542 626614
rect 300986 626058 301222 626294
rect 301306 626058 301542 626294
rect 300986 590378 301222 590614
rect 301306 590378 301542 590614
rect 300986 590058 301222 590294
rect 301306 590058 301542 590294
rect 300986 554378 301222 554614
rect 301306 554378 301542 554614
rect 300986 554058 301222 554294
rect 301306 554058 301542 554294
rect 300986 518378 301222 518614
rect 301306 518378 301542 518614
rect 300986 518058 301222 518294
rect 301306 518058 301542 518294
rect 300986 482378 301222 482614
rect 301306 482378 301542 482614
rect 300986 482058 301222 482294
rect 301306 482058 301542 482294
rect 307826 705562 308062 705798
rect 308146 705562 308382 705798
rect 307826 705242 308062 705478
rect 308146 705242 308382 705478
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 307826 561218 308062 561454
rect 308146 561218 308382 561454
rect 307826 560898 308062 561134
rect 308146 560898 308382 561134
rect 307826 525218 308062 525454
rect 308146 525218 308382 525454
rect 307826 524898 308062 525134
rect 308146 524898 308382 525134
rect 307826 489218 308062 489454
rect 308146 489218 308382 489454
rect 307826 488898 308062 489134
rect 308146 488898 308382 489134
rect 311546 672938 311782 673174
rect 311866 672938 312102 673174
rect 311546 672618 311782 672854
rect 311866 672618 312102 672854
rect 311546 636938 311782 637174
rect 311866 636938 312102 637174
rect 311546 636618 311782 636854
rect 311866 636618 312102 636854
rect 311546 600938 311782 601174
rect 311866 600938 312102 601174
rect 311546 600618 311782 600854
rect 311866 600618 312102 600854
rect 311546 564938 311782 565174
rect 311866 564938 312102 565174
rect 311546 564618 311782 564854
rect 311866 564618 312102 564854
rect 311546 528938 311782 529174
rect 311866 528938 312102 529174
rect 311546 528618 311782 528854
rect 311866 528618 312102 528854
rect 311546 492938 311782 493174
rect 311866 492938 312102 493174
rect 311546 492618 311782 492854
rect 311866 492618 312102 492854
rect 315266 676658 315502 676894
rect 315586 676658 315822 676894
rect 315266 676338 315502 676574
rect 315586 676338 315822 676574
rect 315266 640658 315502 640894
rect 315586 640658 315822 640894
rect 315266 640338 315502 640574
rect 315586 640338 315822 640574
rect 315266 604658 315502 604894
rect 315586 604658 315822 604894
rect 315266 604338 315502 604574
rect 315586 604338 315822 604574
rect 315266 568658 315502 568894
rect 315586 568658 315822 568894
rect 315266 568338 315502 568574
rect 315586 568338 315822 568574
rect 315266 532658 315502 532894
rect 315586 532658 315822 532894
rect 315266 532338 315502 532574
rect 315586 532338 315822 532574
rect 315266 496658 315502 496894
rect 315586 496658 315822 496894
rect 315266 496338 315502 496574
rect 315586 496338 315822 496574
rect 336986 710362 337222 710598
rect 337306 710362 337542 710598
rect 336986 710042 337222 710278
rect 337306 710042 337542 710278
rect 333266 708442 333502 708678
rect 333586 708442 333822 708678
rect 333266 708122 333502 708358
rect 333586 708122 333822 708358
rect 329546 706522 329782 706758
rect 329866 706522 330102 706758
rect 329546 706202 329782 706438
rect 329866 706202 330102 706438
rect 318986 680378 319222 680614
rect 319306 680378 319542 680614
rect 318986 680058 319222 680294
rect 319306 680058 319542 680294
rect 318986 644378 319222 644614
rect 319306 644378 319542 644614
rect 318986 644058 319222 644294
rect 319306 644058 319542 644294
rect 318986 608378 319222 608614
rect 319306 608378 319542 608614
rect 318986 608058 319222 608294
rect 319306 608058 319542 608294
rect 318986 572378 319222 572614
rect 319306 572378 319542 572614
rect 318986 572058 319222 572294
rect 319306 572058 319542 572294
rect 318986 536378 319222 536614
rect 319306 536378 319542 536614
rect 318986 536058 319222 536294
rect 319306 536058 319542 536294
rect 318986 500378 319222 500614
rect 319306 500378 319542 500614
rect 318986 500058 319222 500294
rect 319306 500058 319542 500294
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 325826 543218 326062 543454
rect 326146 543218 326382 543454
rect 325826 542898 326062 543134
rect 326146 542898 326382 543134
rect 325826 507218 326062 507454
rect 326146 507218 326382 507454
rect 325826 506898 326062 507134
rect 326146 506898 326382 507134
rect 329546 690938 329782 691174
rect 329866 690938 330102 691174
rect 329546 690618 329782 690854
rect 329866 690618 330102 690854
rect 329546 654938 329782 655174
rect 329866 654938 330102 655174
rect 329546 654618 329782 654854
rect 329866 654618 330102 654854
rect 329546 618938 329782 619174
rect 329866 618938 330102 619174
rect 329546 618618 329782 618854
rect 329866 618618 330102 618854
rect 329546 582938 329782 583174
rect 329866 582938 330102 583174
rect 329546 582618 329782 582854
rect 329866 582618 330102 582854
rect 329546 546938 329782 547174
rect 329866 546938 330102 547174
rect 329546 546618 329782 546854
rect 329866 546618 330102 546854
rect 329546 510938 329782 511174
rect 329866 510938 330102 511174
rect 329546 510618 329782 510854
rect 329866 510618 330102 510854
rect 333266 694658 333502 694894
rect 333586 694658 333822 694894
rect 333266 694338 333502 694574
rect 333586 694338 333822 694574
rect 333266 658658 333502 658894
rect 333586 658658 333822 658894
rect 333266 658338 333502 658574
rect 333586 658338 333822 658574
rect 333266 622658 333502 622894
rect 333586 622658 333822 622894
rect 333266 622338 333502 622574
rect 333586 622338 333822 622574
rect 333266 586658 333502 586894
rect 333586 586658 333822 586894
rect 333266 586338 333502 586574
rect 333586 586338 333822 586574
rect 333266 550658 333502 550894
rect 333586 550658 333822 550894
rect 333266 550338 333502 550574
rect 333586 550338 333822 550574
rect 333266 514658 333502 514894
rect 333586 514658 333822 514894
rect 333266 514338 333502 514574
rect 333586 514338 333822 514574
rect 354986 711322 355222 711558
rect 355306 711322 355542 711558
rect 354986 711002 355222 711238
rect 355306 711002 355542 711238
rect 351266 709402 351502 709638
rect 351586 709402 351822 709638
rect 351266 709082 351502 709318
rect 351586 709082 351822 709318
rect 347546 707482 347782 707718
rect 347866 707482 348102 707718
rect 347546 707162 347782 707398
rect 347866 707162 348102 707398
rect 336986 698378 337222 698614
rect 337306 698378 337542 698614
rect 336986 698058 337222 698294
rect 337306 698058 337542 698294
rect 336986 662378 337222 662614
rect 337306 662378 337542 662614
rect 336986 662058 337222 662294
rect 337306 662058 337542 662294
rect 336986 626378 337222 626614
rect 337306 626378 337542 626614
rect 336986 626058 337222 626294
rect 337306 626058 337542 626294
rect 336986 590378 337222 590614
rect 337306 590378 337542 590614
rect 336986 590058 337222 590294
rect 337306 590058 337542 590294
rect 336986 554378 337222 554614
rect 337306 554378 337542 554614
rect 336986 554058 337222 554294
rect 337306 554058 337542 554294
rect 336986 518378 337222 518614
rect 337306 518378 337542 518614
rect 336986 518058 337222 518294
rect 337306 518058 337542 518294
rect 336986 482378 337222 482614
rect 337306 482378 337542 482614
rect 336986 482058 337222 482294
rect 337306 482058 337542 482294
rect 343826 705562 344062 705798
rect 344146 705562 344382 705798
rect 343826 705242 344062 705478
rect 344146 705242 344382 705478
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 343826 561218 344062 561454
rect 344146 561218 344382 561454
rect 343826 560898 344062 561134
rect 344146 560898 344382 561134
rect 343826 525218 344062 525454
rect 344146 525218 344382 525454
rect 343826 524898 344062 525134
rect 344146 524898 344382 525134
rect 343826 489218 344062 489454
rect 344146 489218 344382 489454
rect 343826 488898 344062 489134
rect 344146 488898 344382 489134
rect 347546 672938 347782 673174
rect 347866 672938 348102 673174
rect 347546 672618 347782 672854
rect 347866 672618 348102 672854
rect 347546 636938 347782 637174
rect 347866 636938 348102 637174
rect 347546 636618 347782 636854
rect 347866 636618 348102 636854
rect 347546 600938 347782 601174
rect 347866 600938 348102 601174
rect 347546 600618 347782 600854
rect 347866 600618 348102 600854
rect 347546 564938 347782 565174
rect 347866 564938 348102 565174
rect 347546 564618 347782 564854
rect 347866 564618 348102 564854
rect 347546 528938 347782 529174
rect 347866 528938 348102 529174
rect 347546 528618 347782 528854
rect 347866 528618 348102 528854
rect 347546 492938 347782 493174
rect 347866 492938 348102 493174
rect 347546 492618 347782 492854
rect 347866 492618 348102 492854
rect 351266 676658 351502 676894
rect 351586 676658 351822 676894
rect 351266 676338 351502 676574
rect 351586 676338 351822 676574
rect 351266 640658 351502 640894
rect 351586 640658 351822 640894
rect 351266 640338 351502 640574
rect 351586 640338 351822 640574
rect 351266 604658 351502 604894
rect 351586 604658 351822 604894
rect 351266 604338 351502 604574
rect 351586 604338 351822 604574
rect 351266 568658 351502 568894
rect 351586 568658 351822 568894
rect 351266 568338 351502 568574
rect 351586 568338 351822 568574
rect 351266 532658 351502 532894
rect 351586 532658 351822 532894
rect 351266 532338 351502 532574
rect 351586 532338 351822 532574
rect 351266 496658 351502 496894
rect 351586 496658 351822 496894
rect 351266 496338 351502 496574
rect 351586 496338 351822 496574
rect 372986 710362 373222 710598
rect 373306 710362 373542 710598
rect 372986 710042 373222 710278
rect 373306 710042 373542 710278
rect 369266 708442 369502 708678
rect 369586 708442 369822 708678
rect 369266 708122 369502 708358
rect 369586 708122 369822 708358
rect 365546 706522 365782 706758
rect 365866 706522 366102 706758
rect 365546 706202 365782 706438
rect 365866 706202 366102 706438
rect 354986 680378 355222 680614
rect 355306 680378 355542 680614
rect 354986 680058 355222 680294
rect 355306 680058 355542 680294
rect 354986 644378 355222 644614
rect 355306 644378 355542 644614
rect 354986 644058 355222 644294
rect 355306 644058 355542 644294
rect 354986 608378 355222 608614
rect 355306 608378 355542 608614
rect 354986 608058 355222 608294
rect 355306 608058 355542 608294
rect 354986 572378 355222 572614
rect 355306 572378 355542 572614
rect 354986 572058 355222 572294
rect 355306 572058 355542 572294
rect 354986 536378 355222 536614
rect 355306 536378 355542 536614
rect 354986 536058 355222 536294
rect 355306 536058 355542 536294
rect 354986 500378 355222 500614
rect 355306 500378 355542 500614
rect 354986 500058 355222 500294
rect 355306 500058 355542 500294
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 365546 690938 365782 691174
rect 365866 690938 366102 691174
rect 365546 690618 365782 690854
rect 365866 690618 366102 690854
rect 365546 654938 365782 655174
rect 365866 654938 366102 655174
rect 365546 654618 365782 654854
rect 365866 654618 366102 654854
rect 365546 618938 365782 619174
rect 365866 618938 366102 619174
rect 365546 618618 365782 618854
rect 365866 618618 366102 618854
rect 365546 582938 365782 583174
rect 365866 582938 366102 583174
rect 365546 582618 365782 582854
rect 365866 582618 366102 582854
rect 365546 546938 365782 547174
rect 365866 546938 366102 547174
rect 365546 546618 365782 546854
rect 365866 546618 366102 546854
rect 365546 510938 365782 511174
rect 365866 510938 366102 511174
rect 365546 510618 365782 510854
rect 365866 510618 366102 510854
rect 369266 694658 369502 694894
rect 369586 694658 369822 694894
rect 369266 694338 369502 694574
rect 369586 694338 369822 694574
rect 369266 658658 369502 658894
rect 369586 658658 369822 658894
rect 369266 658338 369502 658574
rect 369586 658338 369822 658574
rect 369266 622658 369502 622894
rect 369586 622658 369822 622894
rect 369266 622338 369502 622574
rect 369586 622338 369822 622574
rect 369266 586658 369502 586894
rect 369586 586658 369822 586894
rect 369266 586338 369502 586574
rect 369586 586338 369822 586574
rect 369266 550658 369502 550894
rect 369586 550658 369822 550894
rect 369266 550338 369502 550574
rect 369586 550338 369822 550574
rect 369266 514658 369502 514894
rect 369586 514658 369822 514894
rect 369266 514338 369502 514574
rect 369586 514338 369822 514574
rect 390986 711322 391222 711558
rect 391306 711322 391542 711558
rect 390986 711002 391222 711238
rect 391306 711002 391542 711238
rect 387266 709402 387502 709638
rect 387586 709402 387822 709638
rect 387266 709082 387502 709318
rect 387586 709082 387822 709318
rect 383546 707482 383782 707718
rect 383866 707482 384102 707718
rect 383546 707162 383782 707398
rect 383866 707162 384102 707398
rect 372986 698378 373222 698614
rect 373306 698378 373542 698614
rect 372986 698058 373222 698294
rect 373306 698058 373542 698294
rect 372986 662378 373222 662614
rect 373306 662378 373542 662614
rect 372986 662058 373222 662294
rect 373306 662058 373542 662294
rect 372986 626378 373222 626614
rect 373306 626378 373542 626614
rect 372986 626058 373222 626294
rect 373306 626058 373542 626294
rect 372986 590378 373222 590614
rect 373306 590378 373542 590614
rect 372986 590058 373222 590294
rect 373306 590058 373542 590294
rect 372986 554378 373222 554614
rect 373306 554378 373542 554614
rect 372986 554058 373222 554294
rect 373306 554058 373542 554294
rect 372986 518378 373222 518614
rect 373306 518378 373542 518614
rect 372986 518058 373222 518294
rect 373306 518058 373542 518294
rect 372986 482378 373222 482614
rect 373306 482378 373542 482614
rect 372986 482058 373222 482294
rect 373306 482058 373542 482294
rect 379826 705562 380062 705798
rect 380146 705562 380382 705798
rect 379826 705242 380062 705478
rect 380146 705242 380382 705478
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 379826 561218 380062 561454
rect 380146 561218 380382 561454
rect 379826 560898 380062 561134
rect 380146 560898 380382 561134
rect 379826 525218 380062 525454
rect 380146 525218 380382 525454
rect 379826 524898 380062 525134
rect 380146 524898 380382 525134
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 383546 672938 383782 673174
rect 383866 672938 384102 673174
rect 383546 672618 383782 672854
rect 383866 672618 384102 672854
rect 383546 636938 383782 637174
rect 383866 636938 384102 637174
rect 383546 636618 383782 636854
rect 383866 636618 384102 636854
rect 383546 600938 383782 601174
rect 383866 600938 384102 601174
rect 383546 600618 383782 600854
rect 383866 600618 384102 600854
rect 383546 564938 383782 565174
rect 383866 564938 384102 565174
rect 383546 564618 383782 564854
rect 383866 564618 384102 564854
rect 383546 528938 383782 529174
rect 383866 528938 384102 529174
rect 383546 528618 383782 528854
rect 383866 528618 384102 528854
rect 383546 492938 383782 493174
rect 383866 492938 384102 493174
rect 383546 492618 383782 492854
rect 383866 492618 384102 492854
rect 387266 676658 387502 676894
rect 387586 676658 387822 676894
rect 387266 676338 387502 676574
rect 387586 676338 387822 676574
rect 387266 640658 387502 640894
rect 387586 640658 387822 640894
rect 387266 640338 387502 640574
rect 387586 640338 387822 640574
rect 387266 604658 387502 604894
rect 387586 604658 387822 604894
rect 387266 604338 387502 604574
rect 387586 604338 387822 604574
rect 387266 568658 387502 568894
rect 387586 568658 387822 568894
rect 387266 568338 387502 568574
rect 387586 568338 387822 568574
rect 387266 532658 387502 532894
rect 387586 532658 387822 532894
rect 387266 532338 387502 532574
rect 387586 532338 387822 532574
rect 387266 496658 387502 496894
rect 387586 496658 387822 496894
rect 387266 496338 387502 496574
rect 387586 496338 387822 496574
rect 408986 710362 409222 710598
rect 409306 710362 409542 710598
rect 408986 710042 409222 710278
rect 409306 710042 409542 710278
rect 405266 708442 405502 708678
rect 405586 708442 405822 708678
rect 405266 708122 405502 708358
rect 405586 708122 405822 708358
rect 401546 706522 401782 706758
rect 401866 706522 402102 706758
rect 401546 706202 401782 706438
rect 401866 706202 402102 706438
rect 390986 680378 391222 680614
rect 391306 680378 391542 680614
rect 390986 680058 391222 680294
rect 391306 680058 391542 680294
rect 390986 644378 391222 644614
rect 391306 644378 391542 644614
rect 390986 644058 391222 644294
rect 391306 644058 391542 644294
rect 390986 608378 391222 608614
rect 391306 608378 391542 608614
rect 390986 608058 391222 608294
rect 391306 608058 391542 608294
rect 390986 572378 391222 572614
rect 391306 572378 391542 572614
rect 390986 572058 391222 572294
rect 391306 572058 391542 572294
rect 390986 536378 391222 536614
rect 391306 536378 391542 536614
rect 390986 536058 391222 536294
rect 391306 536058 391542 536294
rect 390986 500378 391222 500614
rect 391306 500378 391542 500614
rect 390986 500058 391222 500294
rect 391306 500058 391542 500294
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 401546 690938 401782 691174
rect 401866 690938 402102 691174
rect 401546 690618 401782 690854
rect 401866 690618 402102 690854
rect 401546 654938 401782 655174
rect 401866 654938 402102 655174
rect 401546 654618 401782 654854
rect 401866 654618 402102 654854
rect 401546 618938 401782 619174
rect 401866 618938 402102 619174
rect 401546 618618 401782 618854
rect 401866 618618 402102 618854
rect 401546 582938 401782 583174
rect 401866 582938 402102 583174
rect 401546 582618 401782 582854
rect 401866 582618 402102 582854
rect 401546 546938 401782 547174
rect 401866 546938 402102 547174
rect 401546 546618 401782 546854
rect 401866 546618 402102 546854
rect 401546 510938 401782 511174
rect 401866 510938 402102 511174
rect 401546 510618 401782 510854
rect 401866 510618 402102 510854
rect 405266 694658 405502 694894
rect 405586 694658 405822 694894
rect 405266 694338 405502 694574
rect 405586 694338 405822 694574
rect 405266 658658 405502 658894
rect 405586 658658 405822 658894
rect 405266 658338 405502 658574
rect 405586 658338 405822 658574
rect 405266 622658 405502 622894
rect 405586 622658 405822 622894
rect 405266 622338 405502 622574
rect 405586 622338 405822 622574
rect 405266 586658 405502 586894
rect 405586 586658 405822 586894
rect 405266 586338 405502 586574
rect 405586 586338 405822 586574
rect 405266 550658 405502 550894
rect 405586 550658 405822 550894
rect 405266 550338 405502 550574
rect 405586 550338 405822 550574
rect 405266 514658 405502 514894
rect 405586 514658 405822 514894
rect 405266 514338 405502 514574
rect 405586 514338 405822 514574
rect 426986 711322 427222 711558
rect 427306 711322 427542 711558
rect 426986 711002 427222 711238
rect 427306 711002 427542 711238
rect 423266 709402 423502 709638
rect 423586 709402 423822 709638
rect 423266 709082 423502 709318
rect 423586 709082 423822 709318
rect 419546 707482 419782 707718
rect 419866 707482 420102 707718
rect 419546 707162 419782 707398
rect 419866 707162 420102 707398
rect 408986 698378 409222 698614
rect 409306 698378 409542 698614
rect 408986 698058 409222 698294
rect 409306 698058 409542 698294
rect 408986 662378 409222 662614
rect 409306 662378 409542 662614
rect 408986 662058 409222 662294
rect 409306 662058 409542 662294
rect 408986 626378 409222 626614
rect 409306 626378 409542 626614
rect 408986 626058 409222 626294
rect 409306 626058 409542 626294
rect 408986 590378 409222 590614
rect 409306 590378 409542 590614
rect 408986 590058 409222 590294
rect 409306 590058 409542 590294
rect 408986 554378 409222 554614
rect 409306 554378 409542 554614
rect 408986 554058 409222 554294
rect 409306 554058 409542 554294
rect 408986 518378 409222 518614
rect 409306 518378 409542 518614
rect 408986 518058 409222 518294
rect 409306 518058 409542 518294
rect 408986 482378 409222 482614
rect 409306 482378 409542 482614
rect 408986 482058 409222 482294
rect 409306 482058 409542 482294
rect 415826 705562 416062 705798
rect 416146 705562 416382 705798
rect 415826 705242 416062 705478
rect 416146 705242 416382 705478
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 415826 561218 416062 561454
rect 416146 561218 416382 561454
rect 415826 560898 416062 561134
rect 416146 560898 416382 561134
rect 415826 525218 416062 525454
rect 416146 525218 416382 525454
rect 415826 524898 416062 525134
rect 416146 524898 416382 525134
rect 415826 489218 416062 489454
rect 416146 489218 416382 489454
rect 415826 488898 416062 489134
rect 416146 488898 416382 489134
rect 419546 672938 419782 673174
rect 419866 672938 420102 673174
rect 419546 672618 419782 672854
rect 419866 672618 420102 672854
rect 419546 636938 419782 637174
rect 419866 636938 420102 637174
rect 419546 636618 419782 636854
rect 419866 636618 420102 636854
rect 419546 600938 419782 601174
rect 419866 600938 420102 601174
rect 419546 600618 419782 600854
rect 419866 600618 420102 600854
rect 419546 564938 419782 565174
rect 419866 564938 420102 565174
rect 419546 564618 419782 564854
rect 419866 564618 420102 564854
rect 419546 528938 419782 529174
rect 419866 528938 420102 529174
rect 419546 528618 419782 528854
rect 419866 528618 420102 528854
rect 419546 492938 419782 493174
rect 419866 492938 420102 493174
rect 419546 492618 419782 492854
rect 419866 492618 420102 492854
rect 423266 676658 423502 676894
rect 423586 676658 423822 676894
rect 423266 676338 423502 676574
rect 423586 676338 423822 676574
rect 423266 640658 423502 640894
rect 423586 640658 423822 640894
rect 423266 640338 423502 640574
rect 423586 640338 423822 640574
rect 423266 604658 423502 604894
rect 423586 604658 423822 604894
rect 423266 604338 423502 604574
rect 423586 604338 423822 604574
rect 423266 568658 423502 568894
rect 423586 568658 423822 568894
rect 423266 568338 423502 568574
rect 423586 568338 423822 568574
rect 423266 532658 423502 532894
rect 423586 532658 423822 532894
rect 423266 532338 423502 532574
rect 423586 532338 423822 532574
rect 423266 496658 423502 496894
rect 423586 496658 423822 496894
rect 423266 496338 423502 496574
rect 423586 496338 423822 496574
rect 444986 710362 445222 710598
rect 445306 710362 445542 710598
rect 444986 710042 445222 710278
rect 445306 710042 445542 710278
rect 441266 708442 441502 708678
rect 441586 708442 441822 708678
rect 441266 708122 441502 708358
rect 441586 708122 441822 708358
rect 437546 706522 437782 706758
rect 437866 706522 438102 706758
rect 437546 706202 437782 706438
rect 437866 706202 438102 706438
rect 426986 680378 427222 680614
rect 427306 680378 427542 680614
rect 426986 680058 427222 680294
rect 427306 680058 427542 680294
rect 426986 644378 427222 644614
rect 427306 644378 427542 644614
rect 426986 644058 427222 644294
rect 427306 644058 427542 644294
rect 426986 608378 427222 608614
rect 427306 608378 427542 608614
rect 426986 608058 427222 608294
rect 427306 608058 427542 608294
rect 426986 572378 427222 572614
rect 427306 572378 427542 572614
rect 426986 572058 427222 572294
rect 427306 572058 427542 572294
rect 426986 536378 427222 536614
rect 427306 536378 427542 536614
rect 426986 536058 427222 536294
rect 427306 536058 427542 536294
rect 426986 500378 427222 500614
rect 427306 500378 427542 500614
rect 426986 500058 427222 500294
rect 427306 500058 427542 500294
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 437546 690938 437782 691174
rect 437866 690938 438102 691174
rect 437546 690618 437782 690854
rect 437866 690618 438102 690854
rect 437546 654938 437782 655174
rect 437866 654938 438102 655174
rect 437546 654618 437782 654854
rect 437866 654618 438102 654854
rect 437546 618938 437782 619174
rect 437866 618938 438102 619174
rect 437546 618618 437782 618854
rect 437866 618618 438102 618854
rect 437546 582938 437782 583174
rect 437866 582938 438102 583174
rect 437546 582618 437782 582854
rect 437866 582618 438102 582854
rect 437546 546938 437782 547174
rect 437866 546938 438102 547174
rect 437546 546618 437782 546854
rect 437866 546618 438102 546854
rect 437546 510938 437782 511174
rect 437866 510938 438102 511174
rect 437546 510618 437782 510854
rect 437866 510618 438102 510854
rect 441266 694658 441502 694894
rect 441586 694658 441822 694894
rect 441266 694338 441502 694574
rect 441586 694338 441822 694574
rect 441266 658658 441502 658894
rect 441586 658658 441822 658894
rect 441266 658338 441502 658574
rect 441586 658338 441822 658574
rect 441266 622658 441502 622894
rect 441586 622658 441822 622894
rect 441266 622338 441502 622574
rect 441586 622338 441822 622574
rect 441266 586658 441502 586894
rect 441586 586658 441822 586894
rect 441266 586338 441502 586574
rect 441586 586338 441822 586574
rect 441266 550658 441502 550894
rect 441586 550658 441822 550894
rect 441266 550338 441502 550574
rect 441586 550338 441822 550574
rect 441266 514658 441502 514894
rect 441586 514658 441822 514894
rect 441266 514338 441502 514574
rect 441586 514338 441822 514574
rect 462986 711322 463222 711558
rect 463306 711322 463542 711558
rect 462986 711002 463222 711238
rect 463306 711002 463542 711238
rect 459266 709402 459502 709638
rect 459586 709402 459822 709638
rect 459266 709082 459502 709318
rect 459586 709082 459822 709318
rect 455546 707482 455782 707718
rect 455866 707482 456102 707718
rect 455546 707162 455782 707398
rect 455866 707162 456102 707398
rect 444986 698378 445222 698614
rect 445306 698378 445542 698614
rect 444986 698058 445222 698294
rect 445306 698058 445542 698294
rect 444986 662378 445222 662614
rect 445306 662378 445542 662614
rect 444986 662058 445222 662294
rect 445306 662058 445542 662294
rect 444986 626378 445222 626614
rect 445306 626378 445542 626614
rect 444986 626058 445222 626294
rect 445306 626058 445542 626294
rect 444986 590378 445222 590614
rect 445306 590378 445542 590614
rect 444986 590058 445222 590294
rect 445306 590058 445542 590294
rect 444986 554378 445222 554614
rect 445306 554378 445542 554614
rect 444986 554058 445222 554294
rect 445306 554058 445542 554294
rect 444986 518378 445222 518614
rect 445306 518378 445542 518614
rect 444986 518058 445222 518294
rect 445306 518058 445542 518294
rect 444986 482378 445222 482614
rect 445306 482378 445542 482614
rect 444986 482058 445222 482294
rect 445306 482058 445542 482294
rect 451826 705562 452062 705798
rect 452146 705562 452382 705798
rect 451826 705242 452062 705478
rect 452146 705242 452382 705478
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 455546 672938 455782 673174
rect 455866 672938 456102 673174
rect 455546 672618 455782 672854
rect 455866 672618 456102 672854
rect 455546 636938 455782 637174
rect 455866 636938 456102 637174
rect 455546 636618 455782 636854
rect 455866 636618 456102 636854
rect 455546 600938 455782 601174
rect 455866 600938 456102 601174
rect 455546 600618 455782 600854
rect 455866 600618 456102 600854
rect 455546 564938 455782 565174
rect 455866 564938 456102 565174
rect 455546 564618 455782 564854
rect 455866 564618 456102 564854
rect 455546 528938 455782 529174
rect 455866 528938 456102 529174
rect 455546 528618 455782 528854
rect 455866 528618 456102 528854
rect 455546 492938 455782 493174
rect 455866 492938 456102 493174
rect 455546 492618 455782 492854
rect 455866 492618 456102 492854
rect 459266 676658 459502 676894
rect 459586 676658 459822 676894
rect 459266 676338 459502 676574
rect 459586 676338 459822 676574
rect 459266 640658 459502 640894
rect 459586 640658 459822 640894
rect 459266 640338 459502 640574
rect 459586 640338 459822 640574
rect 459266 604658 459502 604894
rect 459586 604658 459822 604894
rect 459266 604338 459502 604574
rect 459586 604338 459822 604574
rect 459266 568658 459502 568894
rect 459586 568658 459822 568894
rect 459266 568338 459502 568574
rect 459586 568338 459822 568574
rect 459266 532658 459502 532894
rect 459586 532658 459822 532894
rect 459266 532338 459502 532574
rect 459586 532338 459822 532574
rect 459266 496658 459502 496894
rect 459586 496658 459822 496894
rect 459266 496338 459502 496574
rect 459586 496338 459822 496574
rect 480986 710362 481222 710598
rect 481306 710362 481542 710598
rect 480986 710042 481222 710278
rect 481306 710042 481542 710278
rect 477266 708442 477502 708678
rect 477586 708442 477822 708678
rect 477266 708122 477502 708358
rect 477586 708122 477822 708358
rect 473546 706522 473782 706758
rect 473866 706522 474102 706758
rect 473546 706202 473782 706438
rect 473866 706202 474102 706438
rect 462986 680378 463222 680614
rect 463306 680378 463542 680614
rect 462986 680058 463222 680294
rect 463306 680058 463542 680294
rect 462986 644378 463222 644614
rect 463306 644378 463542 644614
rect 462986 644058 463222 644294
rect 463306 644058 463542 644294
rect 462986 608378 463222 608614
rect 463306 608378 463542 608614
rect 462986 608058 463222 608294
rect 463306 608058 463542 608294
rect 462986 572378 463222 572614
rect 463306 572378 463542 572614
rect 462986 572058 463222 572294
rect 463306 572058 463542 572294
rect 462986 536378 463222 536614
rect 463306 536378 463542 536614
rect 462986 536058 463222 536294
rect 463306 536058 463542 536294
rect 462986 500378 463222 500614
rect 463306 500378 463542 500614
rect 462986 500058 463222 500294
rect 463306 500058 463542 500294
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 473546 690938 473782 691174
rect 473866 690938 474102 691174
rect 473546 690618 473782 690854
rect 473866 690618 474102 690854
rect 473546 654938 473782 655174
rect 473866 654938 474102 655174
rect 473546 654618 473782 654854
rect 473866 654618 474102 654854
rect 473546 618938 473782 619174
rect 473866 618938 474102 619174
rect 473546 618618 473782 618854
rect 473866 618618 474102 618854
rect 473546 582938 473782 583174
rect 473866 582938 474102 583174
rect 473546 582618 473782 582854
rect 473866 582618 474102 582854
rect 473546 546938 473782 547174
rect 473866 546938 474102 547174
rect 473546 546618 473782 546854
rect 473866 546618 474102 546854
rect 473546 510938 473782 511174
rect 473866 510938 474102 511174
rect 473546 510618 473782 510854
rect 473866 510618 474102 510854
rect 477266 694658 477502 694894
rect 477586 694658 477822 694894
rect 477266 694338 477502 694574
rect 477586 694338 477822 694574
rect 477266 658658 477502 658894
rect 477586 658658 477822 658894
rect 477266 658338 477502 658574
rect 477586 658338 477822 658574
rect 477266 622658 477502 622894
rect 477586 622658 477822 622894
rect 477266 622338 477502 622574
rect 477586 622338 477822 622574
rect 477266 586658 477502 586894
rect 477586 586658 477822 586894
rect 477266 586338 477502 586574
rect 477586 586338 477822 586574
rect 477266 550658 477502 550894
rect 477586 550658 477822 550894
rect 477266 550338 477502 550574
rect 477586 550338 477822 550574
rect 477266 514658 477502 514894
rect 477586 514658 477822 514894
rect 477266 514338 477502 514574
rect 477586 514338 477822 514574
rect 498986 711322 499222 711558
rect 499306 711322 499542 711558
rect 498986 711002 499222 711238
rect 499306 711002 499542 711238
rect 495266 709402 495502 709638
rect 495586 709402 495822 709638
rect 495266 709082 495502 709318
rect 495586 709082 495822 709318
rect 491546 707482 491782 707718
rect 491866 707482 492102 707718
rect 491546 707162 491782 707398
rect 491866 707162 492102 707398
rect 480986 698378 481222 698614
rect 481306 698378 481542 698614
rect 480986 698058 481222 698294
rect 481306 698058 481542 698294
rect 480986 662378 481222 662614
rect 481306 662378 481542 662614
rect 480986 662058 481222 662294
rect 481306 662058 481542 662294
rect 480986 626378 481222 626614
rect 481306 626378 481542 626614
rect 480986 626058 481222 626294
rect 481306 626058 481542 626294
rect 480986 590378 481222 590614
rect 481306 590378 481542 590614
rect 480986 590058 481222 590294
rect 481306 590058 481542 590294
rect 480986 554378 481222 554614
rect 481306 554378 481542 554614
rect 480986 554058 481222 554294
rect 481306 554058 481542 554294
rect 480986 518378 481222 518614
rect 481306 518378 481542 518614
rect 480986 518058 481222 518294
rect 481306 518058 481542 518294
rect 480986 482378 481222 482614
rect 481306 482378 481542 482614
rect 480986 482058 481222 482294
rect 481306 482058 481542 482294
rect 487826 705562 488062 705798
rect 488146 705562 488382 705798
rect 487826 705242 488062 705478
rect 488146 705242 488382 705478
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 491546 672938 491782 673174
rect 491866 672938 492102 673174
rect 491546 672618 491782 672854
rect 491866 672618 492102 672854
rect 491546 636938 491782 637174
rect 491866 636938 492102 637174
rect 491546 636618 491782 636854
rect 491866 636618 492102 636854
rect 491546 600938 491782 601174
rect 491866 600938 492102 601174
rect 491546 600618 491782 600854
rect 491866 600618 492102 600854
rect 491546 564938 491782 565174
rect 491866 564938 492102 565174
rect 491546 564618 491782 564854
rect 491866 564618 492102 564854
rect 491546 528938 491782 529174
rect 491866 528938 492102 529174
rect 491546 528618 491782 528854
rect 491866 528618 492102 528854
rect 491546 492938 491782 493174
rect 491866 492938 492102 493174
rect 491546 492618 491782 492854
rect 491866 492618 492102 492854
rect 495266 676658 495502 676894
rect 495586 676658 495822 676894
rect 495266 676338 495502 676574
rect 495586 676338 495822 676574
rect 495266 640658 495502 640894
rect 495586 640658 495822 640894
rect 495266 640338 495502 640574
rect 495586 640338 495822 640574
rect 495266 604658 495502 604894
rect 495586 604658 495822 604894
rect 495266 604338 495502 604574
rect 495586 604338 495822 604574
rect 495266 568658 495502 568894
rect 495586 568658 495822 568894
rect 495266 568338 495502 568574
rect 495586 568338 495822 568574
rect 495266 532658 495502 532894
rect 495586 532658 495822 532894
rect 495266 532338 495502 532574
rect 495586 532338 495822 532574
rect 495266 496658 495502 496894
rect 495586 496658 495822 496894
rect 495266 496338 495502 496574
rect 495586 496338 495822 496574
rect 516986 710362 517222 710598
rect 517306 710362 517542 710598
rect 516986 710042 517222 710278
rect 517306 710042 517542 710278
rect 513266 708442 513502 708678
rect 513586 708442 513822 708678
rect 513266 708122 513502 708358
rect 513586 708122 513822 708358
rect 509546 706522 509782 706758
rect 509866 706522 510102 706758
rect 509546 706202 509782 706438
rect 509866 706202 510102 706438
rect 498986 680378 499222 680614
rect 499306 680378 499542 680614
rect 498986 680058 499222 680294
rect 499306 680058 499542 680294
rect 498986 644378 499222 644614
rect 499306 644378 499542 644614
rect 498986 644058 499222 644294
rect 499306 644058 499542 644294
rect 498986 608378 499222 608614
rect 499306 608378 499542 608614
rect 498986 608058 499222 608294
rect 499306 608058 499542 608294
rect 498986 572378 499222 572614
rect 499306 572378 499542 572614
rect 498986 572058 499222 572294
rect 499306 572058 499542 572294
rect 498986 536378 499222 536614
rect 499306 536378 499542 536614
rect 498986 536058 499222 536294
rect 499306 536058 499542 536294
rect 498986 500378 499222 500614
rect 499306 500378 499542 500614
rect 498986 500058 499222 500294
rect 499306 500058 499542 500294
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 509546 690938 509782 691174
rect 509866 690938 510102 691174
rect 509546 690618 509782 690854
rect 509866 690618 510102 690854
rect 509546 654938 509782 655174
rect 509866 654938 510102 655174
rect 509546 654618 509782 654854
rect 509866 654618 510102 654854
rect 509546 618938 509782 619174
rect 509866 618938 510102 619174
rect 509546 618618 509782 618854
rect 509866 618618 510102 618854
rect 509546 582938 509782 583174
rect 509866 582938 510102 583174
rect 509546 582618 509782 582854
rect 509866 582618 510102 582854
rect 509546 546938 509782 547174
rect 509866 546938 510102 547174
rect 509546 546618 509782 546854
rect 509866 546618 510102 546854
rect 509546 510938 509782 511174
rect 509866 510938 510102 511174
rect 509546 510618 509782 510854
rect 509866 510618 510102 510854
rect 513266 694658 513502 694894
rect 513586 694658 513822 694894
rect 513266 694338 513502 694574
rect 513586 694338 513822 694574
rect 513266 658658 513502 658894
rect 513586 658658 513822 658894
rect 513266 658338 513502 658574
rect 513586 658338 513822 658574
rect 513266 622658 513502 622894
rect 513586 622658 513822 622894
rect 513266 622338 513502 622574
rect 513586 622338 513822 622574
rect 513266 586658 513502 586894
rect 513586 586658 513822 586894
rect 513266 586338 513502 586574
rect 513586 586338 513822 586574
rect 513266 550658 513502 550894
rect 513586 550658 513822 550894
rect 513266 550338 513502 550574
rect 513586 550338 513822 550574
rect 513266 514658 513502 514894
rect 513586 514658 513822 514894
rect 513266 514338 513502 514574
rect 513586 514338 513822 514574
rect 534986 711322 535222 711558
rect 535306 711322 535542 711558
rect 534986 711002 535222 711238
rect 535306 711002 535542 711238
rect 531266 709402 531502 709638
rect 531586 709402 531822 709638
rect 531266 709082 531502 709318
rect 531586 709082 531822 709318
rect 527546 707482 527782 707718
rect 527866 707482 528102 707718
rect 527546 707162 527782 707398
rect 527866 707162 528102 707398
rect 516986 698378 517222 698614
rect 517306 698378 517542 698614
rect 516986 698058 517222 698294
rect 517306 698058 517542 698294
rect 516986 662378 517222 662614
rect 517306 662378 517542 662614
rect 516986 662058 517222 662294
rect 517306 662058 517542 662294
rect 516986 626378 517222 626614
rect 517306 626378 517542 626614
rect 516986 626058 517222 626294
rect 517306 626058 517542 626294
rect 516986 590378 517222 590614
rect 517306 590378 517542 590614
rect 516986 590058 517222 590294
rect 517306 590058 517542 590294
rect 516986 554378 517222 554614
rect 517306 554378 517542 554614
rect 516986 554058 517222 554294
rect 517306 554058 517542 554294
rect 516986 518378 517222 518614
rect 517306 518378 517542 518614
rect 516986 518058 517222 518294
rect 517306 518058 517542 518294
rect 516986 482378 517222 482614
rect 517306 482378 517542 482614
rect 516986 482058 517222 482294
rect 517306 482058 517542 482294
rect 523826 705562 524062 705798
rect 524146 705562 524382 705798
rect 523826 705242 524062 705478
rect 524146 705242 524382 705478
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 527546 672938 527782 673174
rect 527866 672938 528102 673174
rect 527546 672618 527782 672854
rect 527866 672618 528102 672854
rect 527546 636938 527782 637174
rect 527866 636938 528102 637174
rect 527546 636618 527782 636854
rect 527866 636618 528102 636854
rect 527546 600938 527782 601174
rect 527866 600938 528102 601174
rect 527546 600618 527782 600854
rect 527866 600618 528102 600854
rect 527546 564938 527782 565174
rect 527866 564938 528102 565174
rect 527546 564618 527782 564854
rect 527866 564618 528102 564854
rect 527546 528938 527782 529174
rect 527866 528938 528102 529174
rect 527546 528618 527782 528854
rect 527866 528618 528102 528854
rect 527546 492938 527782 493174
rect 527866 492938 528102 493174
rect 527546 492618 527782 492854
rect 527866 492618 528102 492854
rect 531266 676658 531502 676894
rect 531586 676658 531822 676894
rect 531266 676338 531502 676574
rect 531586 676338 531822 676574
rect 531266 640658 531502 640894
rect 531586 640658 531822 640894
rect 531266 640338 531502 640574
rect 531586 640338 531822 640574
rect 531266 604658 531502 604894
rect 531586 604658 531822 604894
rect 531266 604338 531502 604574
rect 531586 604338 531822 604574
rect 531266 568658 531502 568894
rect 531586 568658 531822 568894
rect 531266 568338 531502 568574
rect 531586 568338 531822 568574
rect 531266 532658 531502 532894
rect 531586 532658 531822 532894
rect 531266 532338 531502 532574
rect 531586 532338 531822 532574
rect 531266 496658 531502 496894
rect 531586 496658 531822 496894
rect 531266 496338 531502 496574
rect 531586 496338 531822 496574
rect 552986 710362 553222 710598
rect 553306 710362 553542 710598
rect 552986 710042 553222 710278
rect 553306 710042 553542 710278
rect 549266 708442 549502 708678
rect 549586 708442 549822 708678
rect 549266 708122 549502 708358
rect 549586 708122 549822 708358
rect 545546 706522 545782 706758
rect 545866 706522 546102 706758
rect 545546 706202 545782 706438
rect 545866 706202 546102 706438
rect 534986 680378 535222 680614
rect 535306 680378 535542 680614
rect 534986 680058 535222 680294
rect 535306 680058 535542 680294
rect 534986 644378 535222 644614
rect 535306 644378 535542 644614
rect 534986 644058 535222 644294
rect 535306 644058 535542 644294
rect 534986 608378 535222 608614
rect 535306 608378 535542 608614
rect 534986 608058 535222 608294
rect 535306 608058 535542 608294
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 534986 572378 535222 572614
rect 535306 572378 535542 572614
rect 534986 572058 535222 572294
rect 535306 572058 535542 572294
rect 534986 536378 535222 536614
rect 535306 536378 535542 536614
rect 534986 536058 535222 536294
rect 535306 536058 535542 536294
rect 534986 500378 535222 500614
rect 535306 500378 535542 500614
rect 534986 500058 535222 500294
rect 535306 500058 535542 500294
rect 244250 471218 244486 471454
rect 244250 470898 244486 471134
rect 274970 471218 275206 471454
rect 274970 470898 275206 471134
rect 305690 471218 305926 471454
rect 305690 470898 305926 471134
rect 336410 471218 336646 471454
rect 336410 470898 336646 471134
rect 367130 471218 367366 471454
rect 367130 470898 367366 471134
rect 397850 471218 398086 471454
rect 397850 470898 398086 471134
rect 428570 471218 428806 471454
rect 428570 470898 428806 471134
rect 459290 471218 459526 471454
rect 459290 470898 459526 471134
rect 490010 471218 490246 471454
rect 490010 470898 490246 471134
rect 520730 471218 520966 471454
rect 520730 470898 520966 471134
rect 259610 453218 259846 453454
rect 259610 452898 259846 453134
rect 290330 453218 290566 453454
rect 290330 452898 290566 453134
rect 321050 453218 321286 453454
rect 321050 452898 321286 453134
rect 351770 453218 352006 453454
rect 351770 452898 352006 453134
rect 382490 453218 382726 453454
rect 382490 452898 382726 453134
rect 413210 453218 413446 453454
rect 413210 452898 413446 453134
rect 443930 453218 444166 453454
rect 443930 452898 444166 453134
rect 474650 453218 474886 453454
rect 474650 452898 474886 453134
rect 505370 453218 505606 453454
rect 505370 452898 505606 453134
rect 536090 453218 536326 453454
rect 536090 452898 536326 453134
rect 244250 435218 244486 435454
rect 244250 434898 244486 435134
rect 274970 435218 275206 435454
rect 274970 434898 275206 435134
rect 305690 435218 305926 435454
rect 305690 434898 305926 435134
rect 336410 435218 336646 435454
rect 336410 434898 336646 435134
rect 367130 435218 367366 435454
rect 367130 434898 367366 435134
rect 397850 435218 398086 435454
rect 397850 434898 398086 435134
rect 428570 435218 428806 435454
rect 428570 434898 428806 435134
rect 459290 435218 459526 435454
rect 459290 434898 459526 435134
rect 490010 435218 490246 435454
rect 490010 434898 490246 435134
rect 520730 435218 520966 435454
rect 520730 434898 520966 435134
rect 259610 417218 259846 417454
rect 259610 416898 259846 417134
rect 290330 417218 290566 417454
rect 290330 416898 290566 417134
rect 321050 417218 321286 417454
rect 321050 416898 321286 417134
rect 351770 417218 352006 417454
rect 351770 416898 352006 417134
rect 382490 417218 382726 417454
rect 382490 416898 382726 417134
rect 413210 417218 413446 417454
rect 413210 416898 413446 417134
rect 443930 417218 444166 417454
rect 443930 416898 444166 417134
rect 474650 417218 474886 417454
rect 474650 416898 474886 417134
rect 505370 417218 505606 417454
rect 505370 416898 505606 417134
rect 536090 417218 536326 417454
rect 536090 416898 536326 417134
rect 244250 399218 244486 399454
rect 244250 398898 244486 399134
rect 274970 399218 275206 399454
rect 274970 398898 275206 399134
rect 305690 399218 305926 399454
rect 305690 398898 305926 399134
rect 336410 399218 336646 399454
rect 336410 398898 336646 399134
rect 367130 399218 367366 399454
rect 367130 398898 367366 399134
rect 397850 399218 398086 399454
rect 397850 398898 398086 399134
rect 428570 399218 428806 399454
rect 428570 398898 428806 399134
rect 459290 399218 459526 399454
rect 459290 398898 459526 399134
rect 490010 399218 490246 399454
rect 490010 398898 490246 399134
rect 520730 399218 520966 399454
rect 520730 398898 520966 399134
rect 259610 381218 259846 381454
rect 259610 380898 259846 381134
rect 290330 381218 290566 381454
rect 290330 380898 290566 381134
rect 321050 381218 321286 381454
rect 321050 380898 321286 381134
rect 351770 381218 352006 381454
rect 351770 380898 352006 381134
rect 382490 381218 382726 381454
rect 382490 380898 382726 381134
rect 413210 381218 413446 381454
rect 413210 380898 413446 381134
rect 443930 381218 444166 381454
rect 443930 380898 444166 381134
rect 474650 381218 474886 381454
rect 474650 380898 474886 381134
rect 505370 381218 505606 381454
rect 505370 380898 505606 381134
rect 536090 381218 536326 381454
rect 536090 380898 536326 381134
rect 244250 363218 244486 363454
rect 244250 362898 244486 363134
rect 274970 363218 275206 363454
rect 274970 362898 275206 363134
rect 305690 363218 305926 363454
rect 305690 362898 305926 363134
rect 336410 363218 336646 363454
rect 336410 362898 336646 363134
rect 367130 363218 367366 363454
rect 367130 362898 367366 363134
rect 397850 363218 398086 363454
rect 397850 362898 398086 363134
rect 428570 363218 428806 363454
rect 428570 362898 428806 363134
rect 459290 363218 459526 363454
rect 459290 362898 459526 363134
rect 490010 363218 490246 363454
rect 490010 362898 490246 363134
rect 520730 363218 520966 363454
rect 520730 362898 520966 363134
rect 259610 345218 259846 345454
rect 259610 344898 259846 345134
rect 290330 345218 290566 345454
rect 290330 344898 290566 345134
rect 321050 345218 321286 345454
rect 321050 344898 321286 345134
rect 351770 345218 352006 345454
rect 351770 344898 352006 345134
rect 382490 345218 382726 345454
rect 382490 344898 382726 345134
rect 413210 345218 413446 345454
rect 413210 344898 413446 345134
rect 443930 345218 444166 345454
rect 443930 344898 444166 345134
rect 474650 345218 474886 345454
rect 474650 344898 474886 345134
rect 505370 345218 505606 345454
rect 505370 344898 505606 345134
rect 536090 345218 536326 345454
rect 536090 344898 536326 345134
rect 244250 327218 244486 327454
rect 244250 326898 244486 327134
rect 274970 327218 275206 327454
rect 274970 326898 275206 327134
rect 305690 327218 305926 327454
rect 305690 326898 305926 327134
rect 336410 327218 336646 327454
rect 336410 326898 336646 327134
rect 367130 327218 367366 327454
rect 367130 326898 367366 327134
rect 397850 327218 398086 327454
rect 397850 326898 398086 327134
rect 428570 327218 428806 327454
rect 428570 326898 428806 327134
rect 459290 327218 459526 327454
rect 459290 326898 459526 327134
rect 490010 327218 490246 327454
rect 490010 326898 490246 327134
rect 520730 327218 520966 327454
rect 520730 326898 520966 327134
rect 259610 309218 259846 309454
rect 259610 308898 259846 309134
rect 290330 309218 290566 309454
rect 290330 308898 290566 309134
rect 321050 309218 321286 309454
rect 321050 308898 321286 309134
rect 351770 309218 352006 309454
rect 351770 308898 352006 309134
rect 382490 309218 382726 309454
rect 382490 308898 382726 309134
rect 413210 309218 413446 309454
rect 413210 308898 413446 309134
rect 443930 309218 444166 309454
rect 443930 308898 444166 309134
rect 474650 309218 474886 309454
rect 474650 308898 474886 309134
rect 505370 309218 505606 309454
rect 505370 308898 505606 309134
rect 536090 309218 536326 309454
rect 536090 308898 536326 309134
rect 244250 291218 244486 291454
rect 244250 290898 244486 291134
rect 274970 291218 275206 291454
rect 274970 290898 275206 291134
rect 305690 291218 305926 291454
rect 305690 290898 305926 291134
rect 336410 291218 336646 291454
rect 336410 290898 336646 291134
rect 367130 291218 367366 291454
rect 367130 290898 367366 291134
rect 397850 291218 398086 291454
rect 397850 290898 398086 291134
rect 428570 291218 428806 291454
rect 428570 290898 428806 291134
rect 459290 291218 459526 291454
rect 459290 290898 459526 291134
rect 490010 291218 490246 291454
rect 490010 290898 490246 291134
rect 520730 291218 520966 291454
rect 520730 290898 520966 291134
rect 259610 273218 259846 273454
rect 259610 272898 259846 273134
rect 290330 273218 290566 273454
rect 290330 272898 290566 273134
rect 321050 273218 321286 273454
rect 321050 272898 321286 273134
rect 351770 273218 352006 273454
rect 351770 272898 352006 273134
rect 382490 273218 382726 273454
rect 382490 272898 382726 273134
rect 413210 273218 413446 273454
rect 413210 272898 413446 273134
rect 443930 273218 444166 273454
rect 443930 272898 444166 273134
rect 474650 273218 474886 273454
rect 474650 272898 474886 273134
rect 505370 273218 505606 273454
rect 505370 272898 505606 273134
rect 536090 273218 536326 273454
rect 536090 272898 536326 273134
rect 244250 255218 244486 255454
rect 244250 254898 244486 255134
rect 274970 255218 275206 255454
rect 274970 254898 275206 255134
rect 305690 255218 305926 255454
rect 305690 254898 305926 255134
rect 336410 255218 336646 255454
rect 336410 254898 336646 255134
rect 367130 255218 367366 255454
rect 367130 254898 367366 255134
rect 397850 255218 398086 255454
rect 397850 254898 398086 255134
rect 428570 255218 428806 255454
rect 428570 254898 428806 255134
rect 459290 255218 459526 255454
rect 459290 254898 459526 255134
rect 490010 255218 490246 255454
rect 490010 254898 490246 255134
rect 520730 255218 520966 255454
rect 520730 254898 520966 255134
rect 259610 237218 259846 237454
rect 259610 236898 259846 237134
rect 290330 237218 290566 237454
rect 290330 236898 290566 237134
rect 321050 237218 321286 237454
rect 321050 236898 321286 237134
rect 351770 237218 352006 237454
rect 351770 236898 352006 237134
rect 382490 237218 382726 237454
rect 382490 236898 382726 237134
rect 413210 237218 413446 237454
rect 413210 236898 413446 237134
rect 443930 237218 444166 237454
rect 443930 236898 444166 237134
rect 474650 237218 474886 237454
rect 474650 236898 474886 237134
rect 505370 237218 505606 237454
rect 505370 236898 505606 237134
rect 536090 237218 536326 237454
rect 536090 236898 536326 237134
rect 244250 219218 244486 219454
rect 244250 218898 244486 219134
rect 274970 219218 275206 219454
rect 274970 218898 275206 219134
rect 305690 219218 305926 219454
rect 305690 218898 305926 219134
rect 336410 219218 336646 219454
rect 336410 218898 336646 219134
rect 367130 219218 367366 219454
rect 367130 218898 367366 219134
rect 397850 219218 398086 219454
rect 397850 218898 398086 219134
rect 428570 219218 428806 219454
rect 428570 218898 428806 219134
rect 459290 219218 459526 219454
rect 459290 218898 459526 219134
rect 490010 219218 490246 219454
rect 490010 218898 490246 219134
rect 520730 219218 520966 219454
rect 520730 218898 520966 219134
rect 259610 201218 259846 201454
rect 259610 200898 259846 201134
rect 290330 201218 290566 201454
rect 290330 200898 290566 201134
rect 321050 201218 321286 201454
rect 321050 200898 321286 201134
rect 351770 201218 352006 201454
rect 351770 200898 352006 201134
rect 382490 201218 382726 201454
rect 382490 200898 382726 201134
rect 413210 201218 413446 201454
rect 413210 200898 413446 201134
rect 443930 201218 444166 201454
rect 443930 200898 444166 201134
rect 474650 201218 474886 201454
rect 474650 200898 474886 201134
rect 505370 201218 505606 201454
rect 505370 200898 505606 201134
rect 536090 201218 536326 201454
rect 536090 200898 536326 201134
rect 244250 183218 244486 183454
rect 244250 182898 244486 183134
rect 274970 183218 275206 183454
rect 274970 182898 275206 183134
rect 305690 183218 305926 183454
rect 305690 182898 305926 183134
rect 336410 183218 336646 183454
rect 336410 182898 336646 183134
rect 367130 183218 367366 183454
rect 367130 182898 367366 183134
rect 397850 183218 398086 183454
rect 397850 182898 398086 183134
rect 428570 183218 428806 183454
rect 428570 182898 428806 183134
rect 459290 183218 459526 183454
rect 459290 182898 459526 183134
rect 490010 183218 490246 183454
rect 490010 182898 490246 183134
rect 520730 183218 520966 183454
rect 520730 182898 520966 183134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 545546 690938 545782 691174
rect 545866 690938 546102 691174
rect 545546 690618 545782 690854
rect 545866 690618 546102 690854
rect 545546 654938 545782 655174
rect 545866 654938 546102 655174
rect 545546 654618 545782 654854
rect 545866 654618 546102 654854
rect 545546 618938 545782 619174
rect 545866 618938 546102 619174
rect 545546 618618 545782 618854
rect 545866 618618 546102 618854
rect 545546 582938 545782 583174
rect 545866 582938 546102 583174
rect 545546 582618 545782 582854
rect 545866 582618 546102 582854
rect 545546 546938 545782 547174
rect 545866 546938 546102 547174
rect 545546 546618 545782 546854
rect 545866 546618 546102 546854
rect 545546 510938 545782 511174
rect 545866 510938 546102 511174
rect 545546 510618 545782 510854
rect 545866 510618 546102 510854
rect 545546 474938 545782 475174
rect 545866 474938 546102 475174
rect 545546 474618 545782 474854
rect 545866 474618 546102 474854
rect 545546 438938 545782 439174
rect 545866 438938 546102 439174
rect 545546 438618 545782 438854
rect 545866 438618 546102 438854
rect 545546 402938 545782 403174
rect 545866 402938 546102 403174
rect 545546 402618 545782 402854
rect 545866 402618 546102 402854
rect 545546 366938 545782 367174
rect 545866 366938 546102 367174
rect 545546 366618 545782 366854
rect 545866 366618 546102 366854
rect 545546 330938 545782 331174
rect 545866 330938 546102 331174
rect 545546 330618 545782 330854
rect 545866 330618 546102 330854
rect 545546 294938 545782 295174
rect 545866 294938 546102 295174
rect 545546 294618 545782 294854
rect 545866 294618 546102 294854
rect 545546 258938 545782 259174
rect 545866 258938 546102 259174
rect 545546 258618 545782 258854
rect 545866 258618 546102 258854
rect 545546 222938 545782 223174
rect 545866 222938 546102 223174
rect 545546 222618 545782 222854
rect 545866 222618 546102 222854
rect 545546 186938 545782 187174
rect 545866 186938 546102 187174
rect 545546 186618 545782 186854
rect 545866 186618 546102 186854
rect 235826 165218 236062 165454
rect 236146 165218 236382 165454
rect 235826 164898 236062 165134
rect 236146 164898 236382 165134
rect 235826 129218 236062 129454
rect 236146 129218 236382 129454
rect 235826 128898 236062 129134
rect 236146 128898 236382 129134
rect 235826 93218 236062 93454
rect 236146 93218 236382 93454
rect 235826 92898 236062 93134
rect 236146 92898 236382 93134
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -1542 236062 -1306
rect 236146 -1542 236382 -1306
rect 235826 -1862 236062 -1626
rect 236146 -1862 236382 -1626
rect 239546 168938 239782 169174
rect 239866 168938 240102 169174
rect 239546 168618 239782 168854
rect 239866 168618 240102 168854
rect 239546 132938 239782 133174
rect 239866 132938 240102 133174
rect 239546 132618 239782 132854
rect 239866 132618 240102 132854
rect 239546 96938 239782 97174
rect 239866 96938 240102 97174
rect 239546 96618 239782 96854
rect 239866 96618 240102 96854
rect 239546 60938 239782 61174
rect 239866 60938 240102 61174
rect 239546 60618 239782 60854
rect 239866 60618 240102 60854
rect 239546 24938 239782 25174
rect 239866 24938 240102 25174
rect 239546 24618 239782 24854
rect 239866 24618 240102 24854
rect 239546 -3462 239782 -3226
rect 239866 -3462 240102 -3226
rect 239546 -3782 239782 -3546
rect 239866 -3782 240102 -3546
rect 243266 172658 243502 172894
rect 243586 172658 243822 172894
rect 243266 172338 243502 172574
rect 243586 172338 243822 172574
rect 243266 136658 243502 136894
rect 243586 136658 243822 136894
rect 243266 136338 243502 136574
rect 243586 136338 243822 136574
rect 243266 100658 243502 100894
rect 243586 100658 243822 100894
rect 243266 100338 243502 100574
rect 243586 100338 243822 100574
rect 243266 64658 243502 64894
rect 243586 64658 243822 64894
rect 243266 64338 243502 64574
rect 243586 64338 243822 64574
rect 243266 28658 243502 28894
rect 243586 28658 243822 28894
rect 243266 28338 243502 28574
rect 243586 28338 243822 28574
rect 243266 -5382 243502 -5146
rect 243586 -5382 243822 -5146
rect 243266 -5702 243502 -5466
rect 243586 -5702 243822 -5466
rect 246986 176378 247222 176614
rect 247306 176378 247542 176614
rect 246986 176058 247222 176294
rect 247306 176058 247542 176294
rect 246986 140378 247222 140614
rect 247306 140378 247542 140614
rect 246986 140058 247222 140294
rect 247306 140058 247542 140294
rect 246986 104378 247222 104614
rect 247306 104378 247542 104614
rect 246986 104058 247222 104294
rect 247306 104058 247542 104294
rect 246986 68378 247222 68614
rect 247306 68378 247542 68614
rect 246986 68058 247222 68294
rect 247306 68058 247542 68294
rect 246986 32378 247222 32614
rect 247306 32378 247542 32614
rect 246986 32058 247222 32294
rect 247306 32058 247542 32294
rect 228986 -6342 229222 -6106
rect 229306 -6342 229542 -6106
rect 228986 -6662 229222 -6426
rect 229306 -6662 229542 -6426
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 253826 111218 254062 111454
rect 254146 111218 254382 111454
rect 253826 110898 254062 111134
rect 254146 110898 254382 111134
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 257546 150938 257782 151174
rect 257866 150938 258102 151174
rect 257546 150618 257782 150854
rect 257866 150618 258102 150854
rect 257546 114938 257782 115174
rect 257866 114938 258102 115174
rect 257546 114618 257782 114854
rect 257866 114618 258102 114854
rect 257546 78938 257782 79174
rect 257866 78938 258102 79174
rect 257546 78618 257782 78854
rect 257866 78618 258102 78854
rect 257546 42938 257782 43174
rect 257866 42938 258102 43174
rect 257546 42618 257782 42854
rect 257866 42618 258102 42854
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 257546 -2502 257782 -2266
rect 257866 -2502 258102 -2266
rect 257546 -2822 257782 -2586
rect 257866 -2822 258102 -2586
rect 261266 154658 261502 154894
rect 261586 154658 261822 154894
rect 261266 154338 261502 154574
rect 261586 154338 261822 154574
rect 261266 118658 261502 118894
rect 261586 118658 261822 118894
rect 261266 118338 261502 118574
rect 261586 118338 261822 118574
rect 261266 82658 261502 82894
rect 261586 82658 261822 82894
rect 261266 82338 261502 82574
rect 261586 82338 261822 82574
rect 261266 46658 261502 46894
rect 261586 46658 261822 46894
rect 261266 46338 261502 46574
rect 261586 46338 261822 46574
rect 261266 10658 261502 10894
rect 261586 10658 261822 10894
rect 261266 10338 261502 10574
rect 261586 10338 261822 10574
rect 261266 -4422 261502 -4186
rect 261586 -4422 261822 -4186
rect 261266 -4742 261502 -4506
rect 261586 -4742 261822 -4506
rect 264986 158378 265222 158614
rect 265306 158378 265542 158614
rect 264986 158058 265222 158294
rect 265306 158058 265542 158294
rect 264986 122378 265222 122614
rect 265306 122378 265542 122614
rect 264986 122058 265222 122294
rect 265306 122058 265542 122294
rect 264986 86378 265222 86614
rect 265306 86378 265542 86614
rect 264986 86058 265222 86294
rect 265306 86058 265542 86294
rect 264986 50378 265222 50614
rect 265306 50378 265542 50614
rect 264986 50058 265222 50294
rect 265306 50058 265542 50294
rect 264986 14378 265222 14614
rect 265306 14378 265542 14614
rect 264986 14058 265222 14294
rect 265306 14058 265542 14294
rect 246986 -7302 247222 -7066
rect 247306 -7302 247542 -7066
rect 246986 -7622 247222 -7386
rect 247306 -7622 247542 -7386
rect 271826 165218 272062 165454
rect 272146 165218 272382 165454
rect 271826 164898 272062 165134
rect 272146 164898 272382 165134
rect 271826 129218 272062 129454
rect 272146 129218 272382 129454
rect 271826 128898 272062 129134
rect 272146 128898 272382 129134
rect 271826 93218 272062 93454
rect 272146 93218 272382 93454
rect 271826 92898 272062 93134
rect 272146 92898 272382 93134
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -1542 272062 -1306
rect 272146 -1542 272382 -1306
rect 271826 -1862 272062 -1626
rect 272146 -1862 272382 -1626
rect 275546 168938 275782 169174
rect 275866 168938 276102 169174
rect 275546 168618 275782 168854
rect 275866 168618 276102 168854
rect 275546 132938 275782 133174
rect 275866 132938 276102 133174
rect 275546 132618 275782 132854
rect 275866 132618 276102 132854
rect 275546 96938 275782 97174
rect 275866 96938 276102 97174
rect 275546 96618 275782 96854
rect 275866 96618 276102 96854
rect 275546 60938 275782 61174
rect 275866 60938 276102 61174
rect 275546 60618 275782 60854
rect 275866 60618 276102 60854
rect 275546 24938 275782 25174
rect 275866 24938 276102 25174
rect 275546 24618 275782 24854
rect 275866 24618 276102 24854
rect 275546 -3462 275782 -3226
rect 275866 -3462 276102 -3226
rect 275546 -3782 275782 -3546
rect 275866 -3782 276102 -3546
rect 279266 172658 279502 172894
rect 279586 172658 279822 172894
rect 279266 172338 279502 172574
rect 279586 172338 279822 172574
rect 279266 136658 279502 136894
rect 279586 136658 279822 136894
rect 279266 136338 279502 136574
rect 279586 136338 279822 136574
rect 279266 100658 279502 100894
rect 279586 100658 279822 100894
rect 279266 100338 279502 100574
rect 279586 100338 279822 100574
rect 279266 64658 279502 64894
rect 279586 64658 279822 64894
rect 279266 64338 279502 64574
rect 279586 64338 279822 64574
rect 279266 28658 279502 28894
rect 279586 28658 279822 28894
rect 279266 28338 279502 28574
rect 279586 28338 279822 28574
rect 279266 -5382 279502 -5146
rect 279586 -5382 279822 -5146
rect 279266 -5702 279502 -5466
rect 279586 -5702 279822 -5466
rect 282986 176378 283222 176614
rect 283306 176378 283542 176614
rect 282986 176058 283222 176294
rect 283306 176058 283542 176294
rect 282986 140378 283222 140614
rect 283306 140378 283542 140614
rect 282986 140058 283222 140294
rect 283306 140058 283542 140294
rect 282986 104378 283222 104614
rect 283306 104378 283542 104614
rect 282986 104058 283222 104294
rect 283306 104058 283542 104294
rect 282986 68378 283222 68614
rect 283306 68378 283542 68614
rect 282986 68058 283222 68294
rect 283306 68058 283542 68294
rect 282986 32378 283222 32614
rect 283306 32378 283542 32614
rect 282986 32058 283222 32294
rect 283306 32058 283542 32294
rect 264986 -6342 265222 -6106
rect 265306 -6342 265542 -6106
rect 264986 -6662 265222 -6426
rect 265306 -6662 265542 -6426
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 289826 111218 290062 111454
rect 290146 111218 290382 111454
rect 289826 110898 290062 111134
rect 290146 110898 290382 111134
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 293546 150938 293782 151174
rect 293866 150938 294102 151174
rect 293546 150618 293782 150854
rect 293866 150618 294102 150854
rect 293546 114938 293782 115174
rect 293866 114938 294102 115174
rect 293546 114618 293782 114854
rect 293866 114618 294102 114854
rect 293546 78938 293782 79174
rect 293866 78938 294102 79174
rect 293546 78618 293782 78854
rect 293866 78618 294102 78854
rect 293546 42938 293782 43174
rect 293866 42938 294102 43174
rect 293546 42618 293782 42854
rect 293866 42618 294102 42854
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 293546 -2502 293782 -2266
rect 293866 -2502 294102 -2266
rect 293546 -2822 293782 -2586
rect 293866 -2822 294102 -2586
rect 297266 154658 297502 154894
rect 297586 154658 297822 154894
rect 297266 154338 297502 154574
rect 297586 154338 297822 154574
rect 297266 118658 297502 118894
rect 297586 118658 297822 118894
rect 297266 118338 297502 118574
rect 297586 118338 297822 118574
rect 297266 82658 297502 82894
rect 297586 82658 297822 82894
rect 297266 82338 297502 82574
rect 297586 82338 297822 82574
rect 297266 46658 297502 46894
rect 297586 46658 297822 46894
rect 297266 46338 297502 46574
rect 297586 46338 297822 46574
rect 297266 10658 297502 10894
rect 297586 10658 297822 10894
rect 297266 10338 297502 10574
rect 297586 10338 297822 10574
rect 297266 -4422 297502 -4186
rect 297586 -4422 297822 -4186
rect 297266 -4742 297502 -4506
rect 297586 -4742 297822 -4506
rect 300986 158378 301222 158614
rect 301306 158378 301542 158614
rect 300986 158058 301222 158294
rect 301306 158058 301542 158294
rect 300986 122378 301222 122614
rect 301306 122378 301542 122614
rect 300986 122058 301222 122294
rect 301306 122058 301542 122294
rect 300986 86378 301222 86614
rect 301306 86378 301542 86614
rect 300986 86058 301222 86294
rect 301306 86058 301542 86294
rect 300986 50378 301222 50614
rect 301306 50378 301542 50614
rect 300986 50058 301222 50294
rect 301306 50058 301542 50294
rect 300986 14378 301222 14614
rect 301306 14378 301542 14614
rect 300986 14058 301222 14294
rect 301306 14058 301542 14294
rect 282986 -7302 283222 -7066
rect 283306 -7302 283542 -7066
rect 282986 -7622 283222 -7386
rect 283306 -7622 283542 -7386
rect 307826 165218 308062 165454
rect 308146 165218 308382 165454
rect 307826 164898 308062 165134
rect 308146 164898 308382 165134
rect 307826 129218 308062 129454
rect 308146 129218 308382 129454
rect 307826 128898 308062 129134
rect 308146 128898 308382 129134
rect 307826 93218 308062 93454
rect 308146 93218 308382 93454
rect 307826 92898 308062 93134
rect 308146 92898 308382 93134
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -1542 308062 -1306
rect 308146 -1542 308382 -1306
rect 307826 -1862 308062 -1626
rect 308146 -1862 308382 -1626
rect 311546 168938 311782 169174
rect 311866 168938 312102 169174
rect 311546 168618 311782 168854
rect 311866 168618 312102 168854
rect 311546 132938 311782 133174
rect 311866 132938 312102 133174
rect 311546 132618 311782 132854
rect 311866 132618 312102 132854
rect 311546 96938 311782 97174
rect 311866 96938 312102 97174
rect 311546 96618 311782 96854
rect 311866 96618 312102 96854
rect 311546 60938 311782 61174
rect 311866 60938 312102 61174
rect 311546 60618 311782 60854
rect 311866 60618 312102 60854
rect 311546 24938 311782 25174
rect 311866 24938 312102 25174
rect 311546 24618 311782 24854
rect 311866 24618 312102 24854
rect 311546 -3462 311782 -3226
rect 311866 -3462 312102 -3226
rect 311546 -3782 311782 -3546
rect 311866 -3782 312102 -3546
rect 315266 172658 315502 172894
rect 315586 172658 315822 172894
rect 315266 172338 315502 172574
rect 315586 172338 315822 172574
rect 315266 136658 315502 136894
rect 315586 136658 315822 136894
rect 315266 136338 315502 136574
rect 315586 136338 315822 136574
rect 315266 100658 315502 100894
rect 315586 100658 315822 100894
rect 315266 100338 315502 100574
rect 315586 100338 315822 100574
rect 315266 64658 315502 64894
rect 315586 64658 315822 64894
rect 315266 64338 315502 64574
rect 315586 64338 315822 64574
rect 315266 28658 315502 28894
rect 315586 28658 315822 28894
rect 315266 28338 315502 28574
rect 315586 28338 315822 28574
rect 315266 -5382 315502 -5146
rect 315586 -5382 315822 -5146
rect 315266 -5702 315502 -5466
rect 315586 -5702 315822 -5466
rect 318986 176378 319222 176614
rect 319306 176378 319542 176614
rect 318986 176058 319222 176294
rect 319306 176058 319542 176294
rect 318986 140378 319222 140614
rect 319306 140378 319542 140614
rect 318986 140058 319222 140294
rect 319306 140058 319542 140294
rect 318986 104378 319222 104614
rect 319306 104378 319542 104614
rect 318986 104058 319222 104294
rect 319306 104058 319542 104294
rect 318986 68378 319222 68614
rect 319306 68378 319542 68614
rect 318986 68058 319222 68294
rect 319306 68058 319542 68294
rect 318986 32378 319222 32614
rect 319306 32378 319542 32614
rect 318986 32058 319222 32294
rect 319306 32058 319542 32294
rect 300986 -6342 301222 -6106
rect 301306 -6342 301542 -6106
rect 300986 -6662 301222 -6426
rect 301306 -6662 301542 -6426
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 325826 111218 326062 111454
rect 326146 111218 326382 111454
rect 325826 110898 326062 111134
rect 326146 110898 326382 111134
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 150938 329782 151174
rect 329866 150938 330102 151174
rect 329546 150618 329782 150854
rect 329866 150618 330102 150854
rect 329546 114938 329782 115174
rect 329866 114938 330102 115174
rect 329546 114618 329782 114854
rect 329866 114618 330102 114854
rect 329546 78938 329782 79174
rect 329866 78938 330102 79174
rect 329546 78618 329782 78854
rect 329866 78618 330102 78854
rect 329546 42938 329782 43174
rect 329866 42938 330102 43174
rect 329546 42618 329782 42854
rect 329866 42618 330102 42854
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 329546 -2502 329782 -2266
rect 329866 -2502 330102 -2266
rect 329546 -2822 329782 -2586
rect 329866 -2822 330102 -2586
rect 333266 154658 333502 154894
rect 333586 154658 333822 154894
rect 333266 154338 333502 154574
rect 333586 154338 333822 154574
rect 333266 118658 333502 118894
rect 333586 118658 333822 118894
rect 333266 118338 333502 118574
rect 333586 118338 333822 118574
rect 333266 82658 333502 82894
rect 333586 82658 333822 82894
rect 333266 82338 333502 82574
rect 333586 82338 333822 82574
rect 333266 46658 333502 46894
rect 333586 46658 333822 46894
rect 333266 46338 333502 46574
rect 333586 46338 333822 46574
rect 333266 10658 333502 10894
rect 333586 10658 333822 10894
rect 333266 10338 333502 10574
rect 333586 10338 333822 10574
rect 333266 -4422 333502 -4186
rect 333586 -4422 333822 -4186
rect 333266 -4742 333502 -4506
rect 333586 -4742 333822 -4506
rect 336986 158378 337222 158614
rect 337306 158378 337542 158614
rect 336986 158058 337222 158294
rect 337306 158058 337542 158294
rect 336986 122378 337222 122614
rect 337306 122378 337542 122614
rect 336986 122058 337222 122294
rect 337306 122058 337542 122294
rect 336986 86378 337222 86614
rect 337306 86378 337542 86614
rect 336986 86058 337222 86294
rect 337306 86058 337542 86294
rect 336986 50378 337222 50614
rect 337306 50378 337542 50614
rect 336986 50058 337222 50294
rect 337306 50058 337542 50294
rect 336986 14378 337222 14614
rect 337306 14378 337542 14614
rect 336986 14058 337222 14294
rect 337306 14058 337542 14294
rect 318986 -7302 319222 -7066
rect 319306 -7302 319542 -7066
rect 318986 -7622 319222 -7386
rect 319306 -7622 319542 -7386
rect 343826 165218 344062 165454
rect 344146 165218 344382 165454
rect 343826 164898 344062 165134
rect 344146 164898 344382 165134
rect 343826 129218 344062 129454
rect 344146 129218 344382 129454
rect 343826 128898 344062 129134
rect 344146 128898 344382 129134
rect 343826 93218 344062 93454
rect 344146 93218 344382 93454
rect 343826 92898 344062 93134
rect 344146 92898 344382 93134
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -1542 344062 -1306
rect 344146 -1542 344382 -1306
rect 343826 -1862 344062 -1626
rect 344146 -1862 344382 -1626
rect 347546 168938 347782 169174
rect 347866 168938 348102 169174
rect 347546 168618 347782 168854
rect 347866 168618 348102 168854
rect 347546 132938 347782 133174
rect 347866 132938 348102 133174
rect 347546 132618 347782 132854
rect 347866 132618 348102 132854
rect 347546 96938 347782 97174
rect 347866 96938 348102 97174
rect 347546 96618 347782 96854
rect 347866 96618 348102 96854
rect 347546 60938 347782 61174
rect 347866 60938 348102 61174
rect 347546 60618 347782 60854
rect 347866 60618 348102 60854
rect 347546 24938 347782 25174
rect 347866 24938 348102 25174
rect 347546 24618 347782 24854
rect 347866 24618 348102 24854
rect 347546 -3462 347782 -3226
rect 347866 -3462 348102 -3226
rect 347546 -3782 347782 -3546
rect 347866 -3782 348102 -3546
rect 351266 172658 351502 172894
rect 351586 172658 351822 172894
rect 351266 172338 351502 172574
rect 351586 172338 351822 172574
rect 351266 136658 351502 136894
rect 351586 136658 351822 136894
rect 351266 136338 351502 136574
rect 351586 136338 351822 136574
rect 351266 100658 351502 100894
rect 351586 100658 351822 100894
rect 351266 100338 351502 100574
rect 351586 100338 351822 100574
rect 351266 64658 351502 64894
rect 351586 64658 351822 64894
rect 351266 64338 351502 64574
rect 351586 64338 351822 64574
rect 351266 28658 351502 28894
rect 351586 28658 351822 28894
rect 351266 28338 351502 28574
rect 351586 28338 351822 28574
rect 351266 -5382 351502 -5146
rect 351586 -5382 351822 -5146
rect 351266 -5702 351502 -5466
rect 351586 -5702 351822 -5466
rect 354986 176378 355222 176614
rect 355306 176378 355542 176614
rect 354986 176058 355222 176294
rect 355306 176058 355542 176294
rect 354986 140378 355222 140614
rect 355306 140378 355542 140614
rect 354986 140058 355222 140294
rect 355306 140058 355542 140294
rect 354986 104378 355222 104614
rect 355306 104378 355542 104614
rect 354986 104058 355222 104294
rect 355306 104058 355542 104294
rect 354986 68378 355222 68614
rect 355306 68378 355542 68614
rect 354986 68058 355222 68294
rect 355306 68058 355542 68294
rect 354986 32378 355222 32614
rect 355306 32378 355542 32614
rect 354986 32058 355222 32294
rect 355306 32058 355542 32294
rect 336986 -6342 337222 -6106
rect 337306 -6342 337542 -6106
rect 336986 -6662 337222 -6426
rect 337306 -6662 337542 -6426
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 365546 150938 365782 151174
rect 365866 150938 366102 151174
rect 365546 150618 365782 150854
rect 365866 150618 366102 150854
rect 365546 114938 365782 115174
rect 365866 114938 366102 115174
rect 365546 114618 365782 114854
rect 365866 114618 366102 114854
rect 365546 78938 365782 79174
rect 365866 78938 366102 79174
rect 365546 78618 365782 78854
rect 365866 78618 366102 78854
rect 365546 42938 365782 43174
rect 365866 42938 366102 43174
rect 365546 42618 365782 42854
rect 365866 42618 366102 42854
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 365546 -2502 365782 -2266
rect 365866 -2502 366102 -2266
rect 365546 -2822 365782 -2586
rect 365866 -2822 366102 -2586
rect 369266 154658 369502 154894
rect 369586 154658 369822 154894
rect 369266 154338 369502 154574
rect 369586 154338 369822 154574
rect 369266 118658 369502 118894
rect 369586 118658 369822 118894
rect 369266 118338 369502 118574
rect 369586 118338 369822 118574
rect 369266 82658 369502 82894
rect 369586 82658 369822 82894
rect 369266 82338 369502 82574
rect 369586 82338 369822 82574
rect 369266 46658 369502 46894
rect 369586 46658 369822 46894
rect 369266 46338 369502 46574
rect 369586 46338 369822 46574
rect 369266 10658 369502 10894
rect 369586 10658 369822 10894
rect 369266 10338 369502 10574
rect 369586 10338 369822 10574
rect 369266 -4422 369502 -4186
rect 369586 -4422 369822 -4186
rect 369266 -4742 369502 -4506
rect 369586 -4742 369822 -4506
rect 372986 158378 373222 158614
rect 373306 158378 373542 158614
rect 372986 158058 373222 158294
rect 373306 158058 373542 158294
rect 372986 122378 373222 122614
rect 373306 122378 373542 122614
rect 372986 122058 373222 122294
rect 373306 122058 373542 122294
rect 372986 86378 373222 86614
rect 373306 86378 373542 86614
rect 372986 86058 373222 86294
rect 373306 86058 373542 86294
rect 372986 50378 373222 50614
rect 373306 50378 373542 50614
rect 372986 50058 373222 50294
rect 373306 50058 373542 50294
rect 372986 14378 373222 14614
rect 373306 14378 373542 14614
rect 372986 14058 373222 14294
rect 373306 14058 373542 14294
rect 354986 -7302 355222 -7066
rect 355306 -7302 355542 -7066
rect 354986 -7622 355222 -7386
rect 355306 -7622 355542 -7386
rect 379826 165218 380062 165454
rect 380146 165218 380382 165454
rect 379826 164898 380062 165134
rect 380146 164898 380382 165134
rect 379826 129218 380062 129454
rect 380146 129218 380382 129454
rect 379826 128898 380062 129134
rect 380146 128898 380382 129134
rect 379826 93218 380062 93454
rect 380146 93218 380382 93454
rect 379826 92898 380062 93134
rect 380146 92898 380382 93134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -1542 380062 -1306
rect 380146 -1542 380382 -1306
rect 379826 -1862 380062 -1626
rect 380146 -1862 380382 -1626
rect 383546 168938 383782 169174
rect 383866 168938 384102 169174
rect 383546 168618 383782 168854
rect 383866 168618 384102 168854
rect 383546 132938 383782 133174
rect 383866 132938 384102 133174
rect 383546 132618 383782 132854
rect 383866 132618 384102 132854
rect 383546 96938 383782 97174
rect 383866 96938 384102 97174
rect 383546 96618 383782 96854
rect 383866 96618 384102 96854
rect 383546 60938 383782 61174
rect 383866 60938 384102 61174
rect 383546 60618 383782 60854
rect 383866 60618 384102 60854
rect 383546 24938 383782 25174
rect 383866 24938 384102 25174
rect 383546 24618 383782 24854
rect 383866 24618 384102 24854
rect 383546 -3462 383782 -3226
rect 383866 -3462 384102 -3226
rect 383546 -3782 383782 -3546
rect 383866 -3782 384102 -3546
rect 387266 172658 387502 172894
rect 387586 172658 387822 172894
rect 387266 172338 387502 172574
rect 387586 172338 387822 172574
rect 387266 136658 387502 136894
rect 387586 136658 387822 136894
rect 387266 136338 387502 136574
rect 387586 136338 387822 136574
rect 387266 100658 387502 100894
rect 387586 100658 387822 100894
rect 387266 100338 387502 100574
rect 387586 100338 387822 100574
rect 387266 64658 387502 64894
rect 387586 64658 387822 64894
rect 387266 64338 387502 64574
rect 387586 64338 387822 64574
rect 387266 28658 387502 28894
rect 387586 28658 387822 28894
rect 387266 28338 387502 28574
rect 387586 28338 387822 28574
rect 387266 -5382 387502 -5146
rect 387586 -5382 387822 -5146
rect 387266 -5702 387502 -5466
rect 387586 -5702 387822 -5466
rect 390986 176378 391222 176614
rect 391306 176378 391542 176614
rect 390986 176058 391222 176294
rect 391306 176058 391542 176294
rect 390986 140378 391222 140614
rect 391306 140378 391542 140614
rect 390986 140058 391222 140294
rect 391306 140058 391542 140294
rect 390986 104378 391222 104614
rect 391306 104378 391542 104614
rect 390986 104058 391222 104294
rect 391306 104058 391542 104294
rect 390986 68378 391222 68614
rect 391306 68378 391542 68614
rect 390986 68058 391222 68294
rect 391306 68058 391542 68294
rect 390986 32378 391222 32614
rect 391306 32378 391542 32614
rect 390986 32058 391222 32294
rect 391306 32058 391542 32294
rect 372986 -6342 373222 -6106
rect 373306 -6342 373542 -6106
rect 372986 -6662 373222 -6426
rect 373306 -6662 373542 -6426
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 150938 401782 151174
rect 401866 150938 402102 151174
rect 401546 150618 401782 150854
rect 401866 150618 402102 150854
rect 401546 114938 401782 115174
rect 401866 114938 402102 115174
rect 401546 114618 401782 114854
rect 401866 114618 402102 114854
rect 401546 78938 401782 79174
rect 401866 78938 402102 79174
rect 401546 78618 401782 78854
rect 401866 78618 402102 78854
rect 401546 42938 401782 43174
rect 401866 42938 402102 43174
rect 401546 42618 401782 42854
rect 401866 42618 402102 42854
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -2502 401782 -2266
rect 401866 -2502 402102 -2266
rect 401546 -2822 401782 -2586
rect 401866 -2822 402102 -2586
rect 405266 154658 405502 154894
rect 405586 154658 405822 154894
rect 405266 154338 405502 154574
rect 405586 154338 405822 154574
rect 405266 118658 405502 118894
rect 405586 118658 405822 118894
rect 405266 118338 405502 118574
rect 405586 118338 405822 118574
rect 405266 82658 405502 82894
rect 405586 82658 405822 82894
rect 405266 82338 405502 82574
rect 405586 82338 405822 82574
rect 405266 46658 405502 46894
rect 405586 46658 405822 46894
rect 405266 46338 405502 46574
rect 405586 46338 405822 46574
rect 405266 10658 405502 10894
rect 405586 10658 405822 10894
rect 405266 10338 405502 10574
rect 405586 10338 405822 10574
rect 405266 -4422 405502 -4186
rect 405586 -4422 405822 -4186
rect 405266 -4742 405502 -4506
rect 405586 -4742 405822 -4506
rect 408986 158378 409222 158614
rect 409306 158378 409542 158614
rect 408986 158058 409222 158294
rect 409306 158058 409542 158294
rect 408986 122378 409222 122614
rect 409306 122378 409542 122614
rect 408986 122058 409222 122294
rect 409306 122058 409542 122294
rect 408986 86378 409222 86614
rect 409306 86378 409542 86614
rect 408986 86058 409222 86294
rect 409306 86058 409542 86294
rect 408986 50378 409222 50614
rect 409306 50378 409542 50614
rect 408986 50058 409222 50294
rect 409306 50058 409542 50294
rect 408986 14378 409222 14614
rect 409306 14378 409542 14614
rect 408986 14058 409222 14294
rect 409306 14058 409542 14294
rect 390986 -7302 391222 -7066
rect 391306 -7302 391542 -7066
rect 390986 -7622 391222 -7386
rect 391306 -7622 391542 -7386
rect 415826 165218 416062 165454
rect 416146 165218 416382 165454
rect 415826 164898 416062 165134
rect 416146 164898 416382 165134
rect 415826 129218 416062 129454
rect 416146 129218 416382 129454
rect 415826 128898 416062 129134
rect 416146 128898 416382 129134
rect 415826 93218 416062 93454
rect 416146 93218 416382 93454
rect 415826 92898 416062 93134
rect 416146 92898 416382 93134
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -1542 416062 -1306
rect 416146 -1542 416382 -1306
rect 415826 -1862 416062 -1626
rect 416146 -1862 416382 -1626
rect 419546 168938 419782 169174
rect 419866 168938 420102 169174
rect 419546 168618 419782 168854
rect 419866 168618 420102 168854
rect 419546 132938 419782 133174
rect 419866 132938 420102 133174
rect 419546 132618 419782 132854
rect 419866 132618 420102 132854
rect 419546 96938 419782 97174
rect 419866 96938 420102 97174
rect 419546 96618 419782 96854
rect 419866 96618 420102 96854
rect 419546 60938 419782 61174
rect 419866 60938 420102 61174
rect 419546 60618 419782 60854
rect 419866 60618 420102 60854
rect 419546 24938 419782 25174
rect 419866 24938 420102 25174
rect 419546 24618 419782 24854
rect 419866 24618 420102 24854
rect 419546 -3462 419782 -3226
rect 419866 -3462 420102 -3226
rect 419546 -3782 419782 -3546
rect 419866 -3782 420102 -3546
rect 423266 172658 423502 172894
rect 423586 172658 423822 172894
rect 423266 172338 423502 172574
rect 423586 172338 423822 172574
rect 423266 136658 423502 136894
rect 423586 136658 423822 136894
rect 423266 136338 423502 136574
rect 423586 136338 423822 136574
rect 423266 100658 423502 100894
rect 423586 100658 423822 100894
rect 423266 100338 423502 100574
rect 423586 100338 423822 100574
rect 423266 64658 423502 64894
rect 423586 64658 423822 64894
rect 423266 64338 423502 64574
rect 423586 64338 423822 64574
rect 423266 28658 423502 28894
rect 423586 28658 423822 28894
rect 423266 28338 423502 28574
rect 423586 28338 423822 28574
rect 423266 -5382 423502 -5146
rect 423586 -5382 423822 -5146
rect 423266 -5702 423502 -5466
rect 423586 -5702 423822 -5466
rect 426986 176378 427222 176614
rect 427306 176378 427542 176614
rect 426986 176058 427222 176294
rect 427306 176058 427542 176294
rect 426986 140378 427222 140614
rect 427306 140378 427542 140614
rect 426986 140058 427222 140294
rect 427306 140058 427542 140294
rect 426986 104378 427222 104614
rect 427306 104378 427542 104614
rect 426986 104058 427222 104294
rect 427306 104058 427542 104294
rect 426986 68378 427222 68614
rect 427306 68378 427542 68614
rect 426986 68058 427222 68294
rect 427306 68058 427542 68294
rect 426986 32378 427222 32614
rect 427306 32378 427542 32614
rect 426986 32058 427222 32294
rect 427306 32058 427542 32294
rect 408986 -6342 409222 -6106
rect 409306 -6342 409542 -6106
rect 408986 -6662 409222 -6426
rect 409306 -6662 409542 -6426
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 150938 437782 151174
rect 437866 150938 438102 151174
rect 437546 150618 437782 150854
rect 437866 150618 438102 150854
rect 437546 114938 437782 115174
rect 437866 114938 438102 115174
rect 437546 114618 437782 114854
rect 437866 114618 438102 114854
rect 437546 78938 437782 79174
rect 437866 78938 438102 79174
rect 437546 78618 437782 78854
rect 437866 78618 438102 78854
rect 437546 42938 437782 43174
rect 437866 42938 438102 43174
rect 437546 42618 437782 42854
rect 437866 42618 438102 42854
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 437546 -2502 437782 -2266
rect 437866 -2502 438102 -2266
rect 437546 -2822 437782 -2586
rect 437866 -2822 438102 -2586
rect 441266 154658 441502 154894
rect 441586 154658 441822 154894
rect 441266 154338 441502 154574
rect 441586 154338 441822 154574
rect 441266 118658 441502 118894
rect 441586 118658 441822 118894
rect 441266 118338 441502 118574
rect 441586 118338 441822 118574
rect 441266 82658 441502 82894
rect 441586 82658 441822 82894
rect 441266 82338 441502 82574
rect 441586 82338 441822 82574
rect 441266 46658 441502 46894
rect 441586 46658 441822 46894
rect 441266 46338 441502 46574
rect 441586 46338 441822 46574
rect 441266 10658 441502 10894
rect 441586 10658 441822 10894
rect 441266 10338 441502 10574
rect 441586 10338 441822 10574
rect 441266 -4422 441502 -4186
rect 441586 -4422 441822 -4186
rect 441266 -4742 441502 -4506
rect 441586 -4742 441822 -4506
rect 444986 158378 445222 158614
rect 445306 158378 445542 158614
rect 444986 158058 445222 158294
rect 445306 158058 445542 158294
rect 444986 122378 445222 122614
rect 445306 122378 445542 122614
rect 444986 122058 445222 122294
rect 445306 122058 445542 122294
rect 444986 86378 445222 86614
rect 445306 86378 445542 86614
rect 444986 86058 445222 86294
rect 445306 86058 445542 86294
rect 444986 50378 445222 50614
rect 445306 50378 445542 50614
rect 444986 50058 445222 50294
rect 445306 50058 445542 50294
rect 444986 14378 445222 14614
rect 445306 14378 445542 14614
rect 444986 14058 445222 14294
rect 445306 14058 445542 14294
rect 426986 -7302 427222 -7066
rect 427306 -7302 427542 -7066
rect 426986 -7622 427222 -7386
rect 427306 -7622 427542 -7386
rect 451826 165218 452062 165454
rect 452146 165218 452382 165454
rect 451826 164898 452062 165134
rect 452146 164898 452382 165134
rect 451826 129218 452062 129454
rect 452146 129218 452382 129454
rect 451826 128898 452062 129134
rect 452146 128898 452382 129134
rect 451826 93218 452062 93454
rect 452146 93218 452382 93454
rect 451826 92898 452062 93134
rect 452146 92898 452382 93134
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -1542 452062 -1306
rect 452146 -1542 452382 -1306
rect 451826 -1862 452062 -1626
rect 452146 -1862 452382 -1626
rect 455546 168938 455782 169174
rect 455866 168938 456102 169174
rect 455546 168618 455782 168854
rect 455866 168618 456102 168854
rect 455546 132938 455782 133174
rect 455866 132938 456102 133174
rect 455546 132618 455782 132854
rect 455866 132618 456102 132854
rect 455546 96938 455782 97174
rect 455866 96938 456102 97174
rect 455546 96618 455782 96854
rect 455866 96618 456102 96854
rect 455546 60938 455782 61174
rect 455866 60938 456102 61174
rect 455546 60618 455782 60854
rect 455866 60618 456102 60854
rect 455546 24938 455782 25174
rect 455866 24938 456102 25174
rect 455546 24618 455782 24854
rect 455866 24618 456102 24854
rect 455546 -3462 455782 -3226
rect 455866 -3462 456102 -3226
rect 455546 -3782 455782 -3546
rect 455866 -3782 456102 -3546
rect 459266 172658 459502 172894
rect 459586 172658 459822 172894
rect 459266 172338 459502 172574
rect 459586 172338 459822 172574
rect 459266 136658 459502 136894
rect 459586 136658 459822 136894
rect 459266 136338 459502 136574
rect 459586 136338 459822 136574
rect 459266 100658 459502 100894
rect 459586 100658 459822 100894
rect 459266 100338 459502 100574
rect 459586 100338 459822 100574
rect 459266 64658 459502 64894
rect 459586 64658 459822 64894
rect 459266 64338 459502 64574
rect 459586 64338 459822 64574
rect 459266 28658 459502 28894
rect 459586 28658 459822 28894
rect 459266 28338 459502 28574
rect 459586 28338 459822 28574
rect 459266 -5382 459502 -5146
rect 459586 -5382 459822 -5146
rect 459266 -5702 459502 -5466
rect 459586 -5702 459822 -5466
rect 462986 176378 463222 176614
rect 463306 176378 463542 176614
rect 462986 176058 463222 176294
rect 463306 176058 463542 176294
rect 462986 140378 463222 140614
rect 463306 140378 463542 140614
rect 462986 140058 463222 140294
rect 463306 140058 463542 140294
rect 462986 104378 463222 104614
rect 463306 104378 463542 104614
rect 462986 104058 463222 104294
rect 463306 104058 463542 104294
rect 462986 68378 463222 68614
rect 463306 68378 463542 68614
rect 462986 68058 463222 68294
rect 463306 68058 463542 68294
rect 462986 32378 463222 32614
rect 463306 32378 463542 32614
rect 462986 32058 463222 32294
rect 463306 32058 463542 32294
rect 444986 -6342 445222 -6106
rect 445306 -6342 445542 -6106
rect 444986 -6662 445222 -6426
rect 445306 -6662 445542 -6426
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 150938 473782 151174
rect 473866 150938 474102 151174
rect 473546 150618 473782 150854
rect 473866 150618 474102 150854
rect 473546 114938 473782 115174
rect 473866 114938 474102 115174
rect 473546 114618 473782 114854
rect 473866 114618 474102 114854
rect 473546 78938 473782 79174
rect 473866 78938 474102 79174
rect 473546 78618 473782 78854
rect 473866 78618 474102 78854
rect 473546 42938 473782 43174
rect 473866 42938 474102 43174
rect 473546 42618 473782 42854
rect 473866 42618 474102 42854
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -2502 473782 -2266
rect 473866 -2502 474102 -2266
rect 473546 -2822 473782 -2586
rect 473866 -2822 474102 -2586
rect 477266 154658 477502 154894
rect 477586 154658 477822 154894
rect 477266 154338 477502 154574
rect 477586 154338 477822 154574
rect 477266 118658 477502 118894
rect 477586 118658 477822 118894
rect 477266 118338 477502 118574
rect 477586 118338 477822 118574
rect 477266 82658 477502 82894
rect 477586 82658 477822 82894
rect 477266 82338 477502 82574
rect 477586 82338 477822 82574
rect 477266 46658 477502 46894
rect 477586 46658 477822 46894
rect 477266 46338 477502 46574
rect 477586 46338 477822 46574
rect 477266 10658 477502 10894
rect 477586 10658 477822 10894
rect 477266 10338 477502 10574
rect 477586 10338 477822 10574
rect 477266 -4422 477502 -4186
rect 477586 -4422 477822 -4186
rect 477266 -4742 477502 -4506
rect 477586 -4742 477822 -4506
rect 480986 158378 481222 158614
rect 481306 158378 481542 158614
rect 480986 158058 481222 158294
rect 481306 158058 481542 158294
rect 480986 122378 481222 122614
rect 481306 122378 481542 122614
rect 480986 122058 481222 122294
rect 481306 122058 481542 122294
rect 480986 86378 481222 86614
rect 481306 86378 481542 86614
rect 480986 86058 481222 86294
rect 481306 86058 481542 86294
rect 480986 50378 481222 50614
rect 481306 50378 481542 50614
rect 480986 50058 481222 50294
rect 481306 50058 481542 50294
rect 480986 14378 481222 14614
rect 481306 14378 481542 14614
rect 480986 14058 481222 14294
rect 481306 14058 481542 14294
rect 462986 -7302 463222 -7066
rect 463306 -7302 463542 -7066
rect 462986 -7622 463222 -7386
rect 463306 -7622 463542 -7386
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 487826 129218 488062 129454
rect 488146 129218 488382 129454
rect 487826 128898 488062 129134
rect 488146 128898 488382 129134
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -1542 488062 -1306
rect 488146 -1542 488382 -1306
rect 487826 -1862 488062 -1626
rect 488146 -1862 488382 -1626
rect 491546 168938 491782 169174
rect 491866 168938 492102 169174
rect 491546 168618 491782 168854
rect 491866 168618 492102 168854
rect 491546 132938 491782 133174
rect 491866 132938 492102 133174
rect 491546 132618 491782 132854
rect 491866 132618 492102 132854
rect 491546 96938 491782 97174
rect 491866 96938 492102 97174
rect 491546 96618 491782 96854
rect 491866 96618 492102 96854
rect 491546 60938 491782 61174
rect 491866 60938 492102 61174
rect 491546 60618 491782 60854
rect 491866 60618 492102 60854
rect 491546 24938 491782 25174
rect 491866 24938 492102 25174
rect 491546 24618 491782 24854
rect 491866 24618 492102 24854
rect 491546 -3462 491782 -3226
rect 491866 -3462 492102 -3226
rect 491546 -3782 491782 -3546
rect 491866 -3782 492102 -3546
rect 495266 172658 495502 172894
rect 495586 172658 495822 172894
rect 495266 172338 495502 172574
rect 495586 172338 495822 172574
rect 495266 136658 495502 136894
rect 495586 136658 495822 136894
rect 495266 136338 495502 136574
rect 495586 136338 495822 136574
rect 495266 100658 495502 100894
rect 495586 100658 495822 100894
rect 495266 100338 495502 100574
rect 495586 100338 495822 100574
rect 495266 64658 495502 64894
rect 495586 64658 495822 64894
rect 495266 64338 495502 64574
rect 495586 64338 495822 64574
rect 495266 28658 495502 28894
rect 495586 28658 495822 28894
rect 495266 28338 495502 28574
rect 495586 28338 495822 28574
rect 495266 -5382 495502 -5146
rect 495586 -5382 495822 -5146
rect 495266 -5702 495502 -5466
rect 495586 -5702 495822 -5466
rect 498986 176378 499222 176614
rect 499306 176378 499542 176614
rect 498986 176058 499222 176294
rect 499306 176058 499542 176294
rect 498986 140378 499222 140614
rect 499306 140378 499542 140614
rect 498986 140058 499222 140294
rect 499306 140058 499542 140294
rect 498986 104378 499222 104614
rect 499306 104378 499542 104614
rect 498986 104058 499222 104294
rect 499306 104058 499542 104294
rect 498986 68378 499222 68614
rect 499306 68378 499542 68614
rect 498986 68058 499222 68294
rect 499306 68058 499542 68294
rect 498986 32378 499222 32614
rect 499306 32378 499542 32614
rect 498986 32058 499222 32294
rect 499306 32058 499542 32294
rect 480986 -6342 481222 -6106
rect 481306 -6342 481542 -6106
rect 480986 -6662 481222 -6426
rect 481306 -6662 481542 -6426
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 150938 509782 151174
rect 509866 150938 510102 151174
rect 509546 150618 509782 150854
rect 509866 150618 510102 150854
rect 509546 114938 509782 115174
rect 509866 114938 510102 115174
rect 509546 114618 509782 114854
rect 509866 114618 510102 114854
rect 509546 78938 509782 79174
rect 509866 78938 510102 79174
rect 509546 78618 509782 78854
rect 509866 78618 510102 78854
rect 509546 42938 509782 43174
rect 509866 42938 510102 43174
rect 509546 42618 509782 42854
rect 509866 42618 510102 42854
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -2502 509782 -2266
rect 509866 -2502 510102 -2266
rect 509546 -2822 509782 -2586
rect 509866 -2822 510102 -2586
rect 513266 154658 513502 154894
rect 513586 154658 513822 154894
rect 513266 154338 513502 154574
rect 513586 154338 513822 154574
rect 513266 118658 513502 118894
rect 513586 118658 513822 118894
rect 513266 118338 513502 118574
rect 513586 118338 513822 118574
rect 513266 82658 513502 82894
rect 513586 82658 513822 82894
rect 513266 82338 513502 82574
rect 513586 82338 513822 82574
rect 513266 46658 513502 46894
rect 513586 46658 513822 46894
rect 513266 46338 513502 46574
rect 513586 46338 513822 46574
rect 513266 10658 513502 10894
rect 513586 10658 513822 10894
rect 513266 10338 513502 10574
rect 513586 10338 513822 10574
rect 513266 -4422 513502 -4186
rect 513586 -4422 513822 -4186
rect 513266 -4742 513502 -4506
rect 513586 -4742 513822 -4506
rect 516986 158378 517222 158614
rect 517306 158378 517542 158614
rect 516986 158058 517222 158294
rect 517306 158058 517542 158294
rect 516986 122378 517222 122614
rect 517306 122378 517542 122614
rect 516986 122058 517222 122294
rect 517306 122058 517542 122294
rect 516986 86378 517222 86614
rect 517306 86378 517542 86614
rect 516986 86058 517222 86294
rect 517306 86058 517542 86294
rect 516986 50378 517222 50614
rect 517306 50378 517542 50614
rect 516986 50058 517222 50294
rect 517306 50058 517542 50294
rect 516986 14378 517222 14614
rect 517306 14378 517542 14614
rect 516986 14058 517222 14294
rect 517306 14058 517542 14294
rect 498986 -7302 499222 -7066
rect 499306 -7302 499542 -7066
rect 498986 -7622 499222 -7386
rect 499306 -7622 499542 -7386
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -1542 524062 -1306
rect 524146 -1542 524382 -1306
rect 523826 -1862 524062 -1626
rect 524146 -1862 524382 -1626
rect 527546 168938 527782 169174
rect 527866 168938 528102 169174
rect 527546 168618 527782 168854
rect 527866 168618 528102 168854
rect 527546 132938 527782 133174
rect 527866 132938 528102 133174
rect 527546 132618 527782 132854
rect 527866 132618 528102 132854
rect 527546 96938 527782 97174
rect 527866 96938 528102 97174
rect 527546 96618 527782 96854
rect 527866 96618 528102 96854
rect 527546 60938 527782 61174
rect 527866 60938 528102 61174
rect 527546 60618 527782 60854
rect 527866 60618 528102 60854
rect 527546 24938 527782 25174
rect 527866 24938 528102 25174
rect 527546 24618 527782 24854
rect 527866 24618 528102 24854
rect 527546 -3462 527782 -3226
rect 527866 -3462 528102 -3226
rect 527546 -3782 527782 -3546
rect 527866 -3782 528102 -3546
rect 531266 172658 531502 172894
rect 531586 172658 531822 172894
rect 531266 172338 531502 172574
rect 531586 172338 531822 172574
rect 531266 136658 531502 136894
rect 531586 136658 531822 136894
rect 531266 136338 531502 136574
rect 531586 136338 531822 136574
rect 531266 100658 531502 100894
rect 531586 100658 531822 100894
rect 531266 100338 531502 100574
rect 531586 100338 531822 100574
rect 531266 64658 531502 64894
rect 531586 64658 531822 64894
rect 531266 64338 531502 64574
rect 531586 64338 531822 64574
rect 531266 28658 531502 28894
rect 531586 28658 531822 28894
rect 531266 28338 531502 28574
rect 531586 28338 531822 28574
rect 531266 -5382 531502 -5146
rect 531586 -5382 531822 -5146
rect 531266 -5702 531502 -5466
rect 531586 -5702 531822 -5466
rect 534986 176378 535222 176614
rect 535306 176378 535542 176614
rect 534986 176058 535222 176294
rect 535306 176058 535542 176294
rect 534986 140378 535222 140614
rect 535306 140378 535542 140614
rect 534986 140058 535222 140294
rect 535306 140058 535542 140294
rect 534986 104378 535222 104614
rect 535306 104378 535542 104614
rect 534986 104058 535222 104294
rect 535306 104058 535542 104294
rect 534986 68378 535222 68614
rect 535306 68378 535542 68614
rect 534986 68058 535222 68294
rect 535306 68058 535542 68294
rect 534986 32378 535222 32614
rect 535306 32378 535542 32614
rect 534986 32058 535222 32294
rect 535306 32058 535542 32294
rect 516986 -6342 517222 -6106
rect 517306 -6342 517542 -6106
rect 516986 -6662 517222 -6426
rect 517306 -6662 517542 -6426
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 150938 545782 151174
rect 545866 150938 546102 151174
rect 545546 150618 545782 150854
rect 545866 150618 546102 150854
rect 545546 114938 545782 115174
rect 545866 114938 546102 115174
rect 545546 114618 545782 114854
rect 545866 114618 546102 114854
rect 545546 78938 545782 79174
rect 545866 78938 546102 79174
rect 545546 78618 545782 78854
rect 545866 78618 546102 78854
rect 545546 42938 545782 43174
rect 545866 42938 546102 43174
rect 545546 42618 545782 42854
rect 545866 42618 546102 42854
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -2502 545782 -2266
rect 545866 -2502 546102 -2266
rect 545546 -2822 545782 -2586
rect 545866 -2822 546102 -2586
rect 549266 694658 549502 694894
rect 549586 694658 549822 694894
rect 549266 694338 549502 694574
rect 549586 694338 549822 694574
rect 549266 658658 549502 658894
rect 549586 658658 549822 658894
rect 549266 658338 549502 658574
rect 549586 658338 549822 658574
rect 549266 622658 549502 622894
rect 549586 622658 549822 622894
rect 549266 622338 549502 622574
rect 549586 622338 549822 622574
rect 549266 586658 549502 586894
rect 549586 586658 549822 586894
rect 549266 586338 549502 586574
rect 549586 586338 549822 586574
rect 549266 550658 549502 550894
rect 549586 550658 549822 550894
rect 549266 550338 549502 550574
rect 549586 550338 549822 550574
rect 549266 514658 549502 514894
rect 549586 514658 549822 514894
rect 549266 514338 549502 514574
rect 549586 514338 549822 514574
rect 549266 478658 549502 478894
rect 549586 478658 549822 478894
rect 549266 478338 549502 478574
rect 549586 478338 549822 478574
rect 549266 442658 549502 442894
rect 549586 442658 549822 442894
rect 549266 442338 549502 442574
rect 549586 442338 549822 442574
rect 549266 406658 549502 406894
rect 549586 406658 549822 406894
rect 549266 406338 549502 406574
rect 549586 406338 549822 406574
rect 549266 370658 549502 370894
rect 549586 370658 549822 370894
rect 549266 370338 549502 370574
rect 549586 370338 549822 370574
rect 549266 334658 549502 334894
rect 549586 334658 549822 334894
rect 549266 334338 549502 334574
rect 549586 334338 549822 334574
rect 549266 298658 549502 298894
rect 549586 298658 549822 298894
rect 549266 298338 549502 298574
rect 549586 298338 549822 298574
rect 549266 262658 549502 262894
rect 549586 262658 549822 262894
rect 549266 262338 549502 262574
rect 549586 262338 549822 262574
rect 549266 226658 549502 226894
rect 549586 226658 549822 226894
rect 549266 226338 549502 226574
rect 549586 226338 549822 226574
rect 549266 190658 549502 190894
rect 549586 190658 549822 190894
rect 549266 190338 549502 190574
rect 549586 190338 549822 190574
rect 549266 154658 549502 154894
rect 549586 154658 549822 154894
rect 549266 154338 549502 154574
rect 549586 154338 549822 154574
rect 549266 118658 549502 118894
rect 549586 118658 549822 118894
rect 549266 118338 549502 118574
rect 549586 118338 549822 118574
rect 549266 82658 549502 82894
rect 549586 82658 549822 82894
rect 549266 82338 549502 82574
rect 549586 82338 549822 82574
rect 549266 46658 549502 46894
rect 549586 46658 549822 46894
rect 549266 46338 549502 46574
rect 549586 46338 549822 46574
rect 549266 10658 549502 10894
rect 549586 10658 549822 10894
rect 549266 10338 549502 10574
rect 549586 10338 549822 10574
rect 549266 -4422 549502 -4186
rect 549586 -4422 549822 -4186
rect 549266 -4742 549502 -4506
rect 549586 -4742 549822 -4506
rect 570986 711322 571222 711558
rect 571306 711322 571542 711558
rect 570986 711002 571222 711238
rect 571306 711002 571542 711238
rect 567266 709402 567502 709638
rect 567586 709402 567822 709638
rect 567266 709082 567502 709318
rect 567586 709082 567822 709318
rect 563546 707482 563782 707718
rect 563866 707482 564102 707718
rect 563546 707162 563782 707398
rect 563866 707162 564102 707398
rect 552986 698378 553222 698614
rect 553306 698378 553542 698614
rect 552986 698058 553222 698294
rect 553306 698058 553542 698294
rect 552986 662378 553222 662614
rect 553306 662378 553542 662614
rect 552986 662058 553222 662294
rect 553306 662058 553542 662294
rect 552986 626378 553222 626614
rect 553306 626378 553542 626614
rect 552986 626058 553222 626294
rect 553306 626058 553542 626294
rect 552986 590378 553222 590614
rect 553306 590378 553542 590614
rect 552986 590058 553222 590294
rect 553306 590058 553542 590294
rect 552986 554378 553222 554614
rect 553306 554378 553542 554614
rect 552986 554058 553222 554294
rect 553306 554058 553542 554294
rect 552986 518378 553222 518614
rect 553306 518378 553542 518614
rect 552986 518058 553222 518294
rect 553306 518058 553542 518294
rect 552986 482378 553222 482614
rect 553306 482378 553542 482614
rect 552986 482058 553222 482294
rect 553306 482058 553542 482294
rect 552986 446378 553222 446614
rect 553306 446378 553542 446614
rect 552986 446058 553222 446294
rect 553306 446058 553542 446294
rect 552986 410378 553222 410614
rect 553306 410378 553542 410614
rect 552986 410058 553222 410294
rect 553306 410058 553542 410294
rect 552986 374378 553222 374614
rect 553306 374378 553542 374614
rect 552986 374058 553222 374294
rect 553306 374058 553542 374294
rect 552986 338378 553222 338614
rect 553306 338378 553542 338614
rect 552986 338058 553222 338294
rect 553306 338058 553542 338294
rect 552986 302378 553222 302614
rect 553306 302378 553542 302614
rect 552986 302058 553222 302294
rect 553306 302058 553542 302294
rect 552986 266378 553222 266614
rect 553306 266378 553542 266614
rect 552986 266058 553222 266294
rect 553306 266058 553542 266294
rect 552986 230378 553222 230614
rect 553306 230378 553542 230614
rect 552986 230058 553222 230294
rect 553306 230058 553542 230294
rect 552986 194378 553222 194614
rect 553306 194378 553542 194614
rect 552986 194058 553222 194294
rect 553306 194058 553542 194294
rect 552986 158378 553222 158614
rect 553306 158378 553542 158614
rect 552986 158058 553222 158294
rect 553306 158058 553542 158294
rect 552986 122378 553222 122614
rect 553306 122378 553542 122614
rect 552986 122058 553222 122294
rect 553306 122058 553542 122294
rect 552986 86378 553222 86614
rect 553306 86378 553542 86614
rect 552986 86058 553222 86294
rect 553306 86058 553542 86294
rect 552986 50378 553222 50614
rect 553306 50378 553542 50614
rect 552986 50058 553222 50294
rect 553306 50058 553542 50294
rect 552986 14378 553222 14614
rect 553306 14378 553542 14614
rect 552986 14058 553222 14294
rect 553306 14058 553542 14294
rect 534986 -7302 535222 -7066
rect 535306 -7302 535542 -7066
rect 534986 -7622 535222 -7386
rect 535306 -7622 535542 -7386
rect 559826 705562 560062 705798
rect 560146 705562 560382 705798
rect 559826 705242 560062 705478
rect 560146 705242 560382 705478
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -1542 560062 -1306
rect 560146 -1542 560382 -1306
rect 559826 -1862 560062 -1626
rect 560146 -1862 560382 -1626
rect 563546 672938 563782 673174
rect 563866 672938 564102 673174
rect 563546 672618 563782 672854
rect 563866 672618 564102 672854
rect 563546 636938 563782 637174
rect 563866 636938 564102 637174
rect 563546 636618 563782 636854
rect 563866 636618 564102 636854
rect 563546 600938 563782 601174
rect 563866 600938 564102 601174
rect 563546 600618 563782 600854
rect 563866 600618 564102 600854
rect 563546 564938 563782 565174
rect 563866 564938 564102 565174
rect 563546 564618 563782 564854
rect 563866 564618 564102 564854
rect 563546 528938 563782 529174
rect 563866 528938 564102 529174
rect 563546 528618 563782 528854
rect 563866 528618 564102 528854
rect 563546 492938 563782 493174
rect 563866 492938 564102 493174
rect 563546 492618 563782 492854
rect 563866 492618 564102 492854
rect 563546 456938 563782 457174
rect 563866 456938 564102 457174
rect 563546 456618 563782 456854
rect 563866 456618 564102 456854
rect 563546 420938 563782 421174
rect 563866 420938 564102 421174
rect 563546 420618 563782 420854
rect 563866 420618 564102 420854
rect 563546 384938 563782 385174
rect 563866 384938 564102 385174
rect 563546 384618 563782 384854
rect 563866 384618 564102 384854
rect 563546 348938 563782 349174
rect 563866 348938 564102 349174
rect 563546 348618 563782 348854
rect 563866 348618 564102 348854
rect 563546 312938 563782 313174
rect 563866 312938 564102 313174
rect 563546 312618 563782 312854
rect 563866 312618 564102 312854
rect 563546 276938 563782 277174
rect 563866 276938 564102 277174
rect 563546 276618 563782 276854
rect 563866 276618 564102 276854
rect 563546 240938 563782 241174
rect 563866 240938 564102 241174
rect 563546 240618 563782 240854
rect 563866 240618 564102 240854
rect 563546 204938 563782 205174
rect 563866 204938 564102 205174
rect 563546 204618 563782 204854
rect 563866 204618 564102 204854
rect 563546 168938 563782 169174
rect 563866 168938 564102 169174
rect 563546 168618 563782 168854
rect 563866 168618 564102 168854
rect 563546 132938 563782 133174
rect 563866 132938 564102 133174
rect 563546 132618 563782 132854
rect 563866 132618 564102 132854
rect 563546 96938 563782 97174
rect 563866 96938 564102 97174
rect 563546 96618 563782 96854
rect 563866 96618 564102 96854
rect 563546 60938 563782 61174
rect 563866 60938 564102 61174
rect 563546 60618 563782 60854
rect 563866 60618 564102 60854
rect 563546 24938 563782 25174
rect 563866 24938 564102 25174
rect 563546 24618 563782 24854
rect 563866 24618 564102 24854
rect 563546 -3462 563782 -3226
rect 563866 -3462 564102 -3226
rect 563546 -3782 563782 -3546
rect 563866 -3782 564102 -3546
rect 567266 676658 567502 676894
rect 567586 676658 567822 676894
rect 567266 676338 567502 676574
rect 567586 676338 567822 676574
rect 567266 640658 567502 640894
rect 567586 640658 567822 640894
rect 567266 640338 567502 640574
rect 567586 640338 567822 640574
rect 567266 604658 567502 604894
rect 567586 604658 567822 604894
rect 567266 604338 567502 604574
rect 567586 604338 567822 604574
rect 567266 568658 567502 568894
rect 567586 568658 567822 568894
rect 567266 568338 567502 568574
rect 567586 568338 567822 568574
rect 567266 532658 567502 532894
rect 567586 532658 567822 532894
rect 567266 532338 567502 532574
rect 567586 532338 567822 532574
rect 567266 496658 567502 496894
rect 567586 496658 567822 496894
rect 567266 496338 567502 496574
rect 567586 496338 567822 496574
rect 567266 460658 567502 460894
rect 567586 460658 567822 460894
rect 567266 460338 567502 460574
rect 567586 460338 567822 460574
rect 567266 424658 567502 424894
rect 567586 424658 567822 424894
rect 567266 424338 567502 424574
rect 567586 424338 567822 424574
rect 567266 388658 567502 388894
rect 567586 388658 567822 388894
rect 567266 388338 567502 388574
rect 567586 388338 567822 388574
rect 567266 352658 567502 352894
rect 567586 352658 567822 352894
rect 567266 352338 567502 352574
rect 567586 352338 567822 352574
rect 567266 316658 567502 316894
rect 567586 316658 567822 316894
rect 567266 316338 567502 316574
rect 567586 316338 567822 316574
rect 567266 280658 567502 280894
rect 567586 280658 567822 280894
rect 567266 280338 567502 280574
rect 567586 280338 567822 280574
rect 567266 244658 567502 244894
rect 567586 244658 567822 244894
rect 567266 244338 567502 244574
rect 567586 244338 567822 244574
rect 567266 208658 567502 208894
rect 567586 208658 567822 208894
rect 567266 208338 567502 208574
rect 567586 208338 567822 208574
rect 567266 172658 567502 172894
rect 567586 172658 567822 172894
rect 567266 172338 567502 172574
rect 567586 172338 567822 172574
rect 567266 136658 567502 136894
rect 567586 136658 567822 136894
rect 567266 136338 567502 136574
rect 567586 136338 567822 136574
rect 567266 100658 567502 100894
rect 567586 100658 567822 100894
rect 567266 100338 567502 100574
rect 567586 100338 567822 100574
rect 567266 64658 567502 64894
rect 567586 64658 567822 64894
rect 567266 64338 567502 64574
rect 567586 64338 567822 64574
rect 567266 28658 567502 28894
rect 567586 28658 567822 28894
rect 567266 28338 567502 28574
rect 567586 28338 567822 28574
rect 567266 -5382 567502 -5146
rect 567586 -5382 567822 -5146
rect 567266 -5702 567502 -5466
rect 567586 -5702 567822 -5466
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 581546 706522 581782 706758
rect 581866 706522 582102 706758
rect 581546 706202 581782 706438
rect 581866 706202 582102 706438
rect 570986 680378 571222 680614
rect 571306 680378 571542 680614
rect 570986 680058 571222 680294
rect 571306 680058 571542 680294
rect 570986 644378 571222 644614
rect 571306 644378 571542 644614
rect 570986 644058 571222 644294
rect 571306 644058 571542 644294
rect 570986 608378 571222 608614
rect 571306 608378 571542 608614
rect 570986 608058 571222 608294
rect 571306 608058 571542 608294
rect 570986 572378 571222 572614
rect 571306 572378 571542 572614
rect 570986 572058 571222 572294
rect 571306 572058 571542 572294
rect 570986 536378 571222 536614
rect 571306 536378 571542 536614
rect 570986 536058 571222 536294
rect 571306 536058 571542 536294
rect 570986 500378 571222 500614
rect 571306 500378 571542 500614
rect 570986 500058 571222 500294
rect 571306 500058 571542 500294
rect 570986 464378 571222 464614
rect 571306 464378 571542 464614
rect 570986 464058 571222 464294
rect 571306 464058 571542 464294
rect 570986 428378 571222 428614
rect 571306 428378 571542 428614
rect 570986 428058 571222 428294
rect 571306 428058 571542 428294
rect 570986 392378 571222 392614
rect 571306 392378 571542 392614
rect 570986 392058 571222 392294
rect 571306 392058 571542 392294
rect 570986 356378 571222 356614
rect 571306 356378 571542 356614
rect 570986 356058 571222 356294
rect 571306 356058 571542 356294
rect 570986 320378 571222 320614
rect 571306 320378 571542 320614
rect 570986 320058 571222 320294
rect 571306 320058 571542 320294
rect 570986 284378 571222 284614
rect 571306 284378 571542 284614
rect 570986 284058 571222 284294
rect 571306 284058 571542 284294
rect 570986 248378 571222 248614
rect 571306 248378 571542 248614
rect 570986 248058 571222 248294
rect 571306 248058 571542 248294
rect 570986 212378 571222 212614
rect 571306 212378 571542 212614
rect 570986 212058 571222 212294
rect 571306 212058 571542 212294
rect 570986 176378 571222 176614
rect 571306 176378 571542 176614
rect 570986 176058 571222 176294
rect 571306 176058 571542 176294
rect 570986 140378 571222 140614
rect 571306 140378 571542 140614
rect 570986 140058 571222 140294
rect 571306 140058 571542 140294
rect 570986 104378 571222 104614
rect 571306 104378 571542 104614
rect 570986 104058 571222 104294
rect 571306 104058 571542 104294
rect 570986 68378 571222 68614
rect 571306 68378 571542 68614
rect 570986 68058 571222 68294
rect 571306 68058 571542 68294
rect 570986 32378 571222 32614
rect 571306 32378 571542 32614
rect 570986 32058 571222 32294
rect 571306 32058 571542 32294
rect 552986 -6342 553222 -6106
rect 553306 -6342 553542 -6106
rect 552986 -6662 553222 -6426
rect 553306 -6662 553542 -6426
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 669218 586538 669454
rect 586622 669218 586858 669454
rect 586302 668898 586538 669134
rect 586622 668898 586858 669134
rect 586302 633218 586538 633454
rect 586622 633218 586858 633454
rect 586302 632898 586538 633134
rect 586622 632898 586858 633134
rect 586302 597218 586538 597454
rect 586622 597218 586858 597454
rect 586302 596898 586538 597134
rect 586622 596898 586858 597134
rect 586302 561218 586538 561454
rect 586622 561218 586858 561454
rect 586302 560898 586538 561134
rect 586622 560898 586858 561134
rect 586302 525218 586538 525454
rect 586622 525218 586858 525454
rect 586302 524898 586538 525134
rect 586622 524898 586858 525134
rect 586302 489218 586538 489454
rect 586622 489218 586858 489454
rect 586302 488898 586538 489134
rect 586622 488898 586858 489134
rect 586302 453218 586538 453454
rect 586622 453218 586858 453454
rect 586302 452898 586538 453134
rect 586622 452898 586858 453134
rect 586302 417218 586538 417454
rect 586622 417218 586858 417454
rect 586302 416898 586538 417134
rect 586622 416898 586858 417134
rect 586302 381218 586538 381454
rect 586622 381218 586858 381454
rect 586302 380898 586538 381134
rect 586622 380898 586858 381134
rect 586302 345218 586538 345454
rect 586622 345218 586858 345454
rect 586302 344898 586538 345134
rect 586622 344898 586858 345134
rect 586302 309218 586538 309454
rect 586622 309218 586858 309454
rect 586302 308898 586538 309134
rect 586622 308898 586858 309134
rect 586302 273218 586538 273454
rect 586622 273218 586858 273454
rect 586302 272898 586538 273134
rect 586622 272898 586858 273134
rect 586302 237218 586538 237454
rect 586622 237218 586858 237454
rect 586302 236898 586538 237134
rect 586622 236898 586858 237134
rect 586302 201218 586538 201454
rect 586622 201218 586858 201454
rect 586302 200898 586538 201134
rect 586622 200898 586858 201134
rect 586302 165218 586538 165454
rect 586622 165218 586858 165454
rect 586302 164898 586538 165134
rect 586622 164898 586858 165134
rect 586302 129218 586538 129454
rect 586622 129218 586858 129454
rect 586302 128898 586538 129134
rect 586622 128898 586858 129134
rect 586302 93218 586538 93454
rect 586622 93218 586858 93454
rect 586302 92898 586538 93134
rect 586622 92898 586858 93134
rect 586302 57218 586538 57454
rect 586622 57218 586858 57454
rect 586302 56898 586538 57134
rect 586622 56898 586858 57134
rect 586302 21218 586538 21454
rect 586622 21218 586858 21454
rect 586302 20898 586538 21134
rect 586622 20898 586858 21134
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 690938 587498 691174
rect 587582 690938 587818 691174
rect 587262 690618 587498 690854
rect 587582 690618 587818 690854
rect 587262 654938 587498 655174
rect 587582 654938 587818 655174
rect 587262 654618 587498 654854
rect 587582 654618 587818 654854
rect 587262 618938 587498 619174
rect 587582 618938 587818 619174
rect 587262 618618 587498 618854
rect 587582 618618 587818 618854
rect 587262 582938 587498 583174
rect 587582 582938 587818 583174
rect 587262 582618 587498 582854
rect 587582 582618 587818 582854
rect 587262 546938 587498 547174
rect 587582 546938 587818 547174
rect 587262 546618 587498 546854
rect 587582 546618 587818 546854
rect 587262 510938 587498 511174
rect 587582 510938 587818 511174
rect 587262 510618 587498 510854
rect 587582 510618 587818 510854
rect 587262 474938 587498 475174
rect 587582 474938 587818 475174
rect 587262 474618 587498 474854
rect 587582 474618 587818 474854
rect 587262 438938 587498 439174
rect 587582 438938 587818 439174
rect 587262 438618 587498 438854
rect 587582 438618 587818 438854
rect 587262 402938 587498 403174
rect 587582 402938 587818 403174
rect 587262 402618 587498 402854
rect 587582 402618 587818 402854
rect 587262 366938 587498 367174
rect 587582 366938 587818 367174
rect 587262 366618 587498 366854
rect 587582 366618 587818 366854
rect 587262 330938 587498 331174
rect 587582 330938 587818 331174
rect 587262 330618 587498 330854
rect 587582 330618 587818 330854
rect 587262 294938 587498 295174
rect 587582 294938 587818 295174
rect 587262 294618 587498 294854
rect 587582 294618 587818 294854
rect 587262 258938 587498 259174
rect 587582 258938 587818 259174
rect 587262 258618 587498 258854
rect 587582 258618 587818 258854
rect 587262 222938 587498 223174
rect 587582 222938 587818 223174
rect 587262 222618 587498 222854
rect 587582 222618 587818 222854
rect 587262 186938 587498 187174
rect 587582 186938 587818 187174
rect 587262 186618 587498 186854
rect 587582 186618 587818 186854
rect 587262 150938 587498 151174
rect 587582 150938 587818 151174
rect 587262 150618 587498 150854
rect 587582 150618 587818 150854
rect 587262 114938 587498 115174
rect 587582 114938 587818 115174
rect 587262 114618 587498 114854
rect 587582 114618 587818 114854
rect 587262 78938 587498 79174
rect 587582 78938 587818 79174
rect 587262 78618 587498 78854
rect 587582 78618 587818 78854
rect 587262 42938 587498 43174
rect 587582 42938 587818 43174
rect 587262 42618 587498 42854
rect 587582 42618 587818 42854
rect 587262 6938 587498 7174
rect 587582 6938 587818 7174
rect 587262 6618 587498 6854
rect 587582 6618 587818 6854
rect 581546 -2502 581782 -2266
rect 581866 -2502 582102 -2266
rect 581546 -2822 581782 -2586
rect 581866 -2822 582102 -2586
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 672938 588458 673174
rect 588542 672938 588778 673174
rect 588222 672618 588458 672854
rect 588542 672618 588778 672854
rect 588222 636938 588458 637174
rect 588542 636938 588778 637174
rect 588222 636618 588458 636854
rect 588542 636618 588778 636854
rect 588222 600938 588458 601174
rect 588542 600938 588778 601174
rect 588222 600618 588458 600854
rect 588542 600618 588778 600854
rect 588222 564938 588458 565174
rect 588542 564938 588778 565174
rect 588222 564618 588458 564854
rect 588542 564618 588778 564854
rect 588222 528938 588458 529174
rect 588542 528938 588778 529174
rect 588222 528618 588458 528854
rect 588542 528618 588778 528854
rect 588222 492938 588458 493174
rect 588542 492938 588778 493174
rect 588222 492618 588458 492854
rect 588542 492618 588778 492854
rect 588222 456938 588458 457174
rect 588542 456938 588778 457174
rect 588222 456618 588458 456854
rect 588542 456618 588778 456854
rect 588222 420938 588458 421174
rect 588542 420938 588778 421174
rect 588222 420618 588458 420854
rect 588542 420618 588778 420854
rect 588222 384938 588458 385174
rect 588542 384938 588778 385174
rect 588222 384618 588458 384854
rect 588542 384618 588778 384854
rect 588222 348938 588458 349174
rect 588542 348938 588778 349174
rect 588222 348618 588458 348854
rect 588542 348618 588778 348854
rect 588222 312938 588458 313174
rect 588542 312938 588778 313174
rect 588222 312618 588458 312854
rect 588542 312618 588778 312854
rect 588222 276938 588458 277174
rect 588542 276938 588778 277174
rect 588222 276618 588458 276854
rect 588542 276618 588778 276854
rect 588222 240938 588458 241174
rect 588542 240938 588778 241174
rect 588222 240618 588458 240854
rect 588542 240618 588778 240854
rect 588222 204938 588458 205174
rect 588542 204938 588778 205174
rect 588222 204618 588458 204854
rect 588542 204618 588778 204854
rect 588222 168938 588458 169174
rect 588542 168938 588778 169174
rect 588222 168618 588458 168854
rect 588542 168618 588778 168854
rect 588222 132938 588458 133174
rect 588542 132938 588778 133174
rect 588222 132618 588458 132854
rect 588542 132618 588778 132854
rect 588222 96938 588458 97174
rect 588542 96938 588778 97174
rect 588222 96618 588458 96854
rect 588542 96618 588778 96854
rect 588222 60938 588458 61174
rect 588542 60938 588778 61174
rect 588222 60618 588458 60854
rect 588542 60618 588778 60854
rect 588222 24938 588458 25174
rect 588542 24938 588778 25174
rect 588222 24618 588458 24854
rect 588542 24618 588778 24854
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 694658 589418 694894
rect 589502 694658 589738 694894
rect 589182 694338 589418 694574
rect 589502 694338 589738 694574
rect 589182 658658 589418 658894
rect 589502 658658 589738 658894
rect 589182 658338 589418 658574
rect 589502 658338 589738 658574
rect 589182 622658 589418 622894
rect 589502 622658 589738 622894
rect 589182 622338 589418 622574
rect 589502 622338 589738 622574
rect 589182 586658 589418 586894
rect 589502 586658 589738 586894
rect 589182 586338 589418 586574
rect 589502 586338 589738 586574
rect 589182 550658 589418 550894
rect 589502 550658 589738 550894
rect 589182 550338 589418 550574
rect 589502 550338 589738 550574
rect 589182 514658 589418 514894
rect 589502 514658 589738 514894
rect 589182 514338 589418 514574
rect 589502 514338 589738 514574
rect 589182 478658 589418 478894
rect 589502 478658 589738 478894
rect 589182 478338 589418 478574
rect 589502 478338 589738 478574
rect 589182 442658 589418 442894
rect 589502 442658 589738 442894
rect 589182 442338 589418 442574
rect 589502 442338 589738 442574
rect 589182 406658 589418 406894
rect 589502 406658 589738 406894
rect 589182 406338 589418 406574
rect 589502 406338 589738 406574
rect 589182 370658 589418 370894
rect 589502 370658 589738 370894
rect 589182 370338 589418 370574
rect 589502 370338 589738 370574
rect 589182 334658 589418 334894
rect 589502 334658 589738 334894
rect 589182 334338 589418 334574
rect 589502 334338 589738 334574
rect 589182 298658 589418 298894
rect 589502 298658 589738 298894
rect 589182 298338 589418 298574
rect 589502 298338 589738 298574
rect 589182 262658 589418 262894
rect 589502 262658 589738 262894
rect 589182 262338 589418 262574
rect 589502 262338 589738 262574
rect 589182 226658 589418 226894
rect 589502 226658 589738 226894
rect 589182 226338 589418 226574
rect 589502 226338 589738 226574
rect 589182 190658 589418 190894
rect 589502 190658 589738 190894
rect 589182 190338 589418 190574
rect 589502 190338 589738 190574
rect 589182 154658 589418 154894
rect 589502 154658 589738 154894
rect 589182 154338 589418 154574
rect 589502 154338 589738 154574
rect 589182 118658 589418 118894
rect 589502 118658 589738 118894
rect 589182 118338 589418 118574
rect 589502 118338 589738 118574
rect 589182 82658 589418 82894
rect 589502 82658 589738 82894
rect 589182 82338 589418 82574
rect 589502 82338 589738 82574
rect 589182 46658 589418 46894
rect 589502 46658 589738 46894
rect 589182 46338 589418 46574
rect 589502 46338 589738 46574
rect 589182 10658 589418 10894
rect 589502 10658 589738 10894
rect 589182 10338 589418 10574
rect 589502 10338 589738 10574
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 676658 590378 676894
rect 590462 676658 590698 676894
rect 590142 676338 590378 676574
rect 590462 676338 590698 676574
rect 590142 640658 590378 640894
rect 590462 640658 590698 640894
rect 590142 640338 590378 640574
rect 590462 640338 590698 640574
rect 590142 604658 590378 604894
rect 590462 604658 590698 604894
rect 590142 604338 590378 604574
rect 590462 604338 590698 604574
rect 590142 568658 590378 568894
rect 590462 568658 590698 568894
rect 590142 568338 590378 568574
rect 590462 568338 590698 568574
rect 590142 532658 590378 532894
rect 590462 532658 590698 532894
rect 590142 532338 590378 532574
rect 590462 532338 590698 532574
rect 590142 496658 590378 496894
rect 590462 496658 590698 496894
rect 590142 496338 590378 496574
rect 590462 496338 590698 496574
rect 590142 460658 590378 460894
rect 590462 460658 590698 460894
rect 590142 460338 590378 460574
rect 590462 460338 590698 460574
rect 590142 424658 590378 424894
rect 590462 424658 590698 424894
rect 590142 424338 590378 424574
rect 590462 424338 590698 424574
rect 590142 388658 590378 388894
rect 590462 388658 590698 388894
rect 590142 388338 590378 388574
rect 590462 388338 590698 388574
rect 590142 352658 590378 352894
rect 590462 352658 590698 352894
rect 590142 352338 590378 352574
rect 590462 352338 590698 352574
rect 590142 316658 590378 316894
rect 590462 316658 590698 316894
rect 590142 316338 590378 316574
rect 590462 316338 590698 316574
rect 590142 280658 590378 280894
rect 590462 280658 590698 280894
rect 590142 280338 590378 280574
rect 590462 280338 590698 280574
rect 590142 244658 590378 244894
rect 590462 244658 590698 244894
rect 590142 244338 590378 244574
rect 590462 244338 590698 244574
rect 590142 208658 590378 208894
rect 590462 208658 590698 208894
rect 590142 208338 590378 208574
rect 590462 208338 590698 208574
rect 590142 172658 590378 172894
rect 590462 172658 590698 172894
rect 590142 172338 590378 172574
rect 590462 172338 590698 172574
rect 590142 136658 590378 136894
rect 590462 136658 590698 136894
rect 590142 136338 590378 136574
rect 590462 136338 590698 136574
rect 590142 100658 590378 100894
rect 590462 100658 590698 100894
rect 590142 100338 590378 100574
rect 590462 100338 590698 100574
rect 590142 64658 590378 64894
rect 590462 64658 590698 64894
rect 590142 64338 590378 64574
rect 590462 64338 590698 64574
rect 590142 28658 590378 28894
rect 590462 28658 590698 28894
rect 590142 28338 590378 28574
rect 590462 28338 590698 28574
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 698378 591338 698614
rect 591422 698378 591658 698614
rect 591102 698058 591338 698294
rect 591422 698058 591658 698294
rect 591102 662378 591338 662614
rect 591422 662378 591658 662614
rect 591102 662058 591338 662294
rect 591422 662058 591658 662294
rect 591102 626378 591338 626614
rect 591422 626378 591658 626614
rect 591102 626058 591338 626294
rect 591422 626058 591658 626294
rect 591102 590378 591338 590614
rect 591422 590378 591658 590614
rect 591102 590058 591338 590294
rect 591422 590058 591658 590294
rect 591102 554378 591338 554614
rect 591422 554378 591658 554614
rect 591102 554058 591338 554294
rect 591422 554058 591658 554294
rect 591102 518378 591338 518614
rect 591422 518378 591658 518614
rect 591102 518058 591338 518294
rect 591422 518058 591658 518294
rect 591102 482378 591338 482614
rect 591422 482378 591658 482614
rect 591102 482058 591338 482294
rect 591422 482058 591658 482294
rect 591102 446378 591338 446614
rect 591422 446378 591658 446614
rect 591102 446058 591338 446294
rect 591422 446058 591658 446294
rect 591102 410378 591338 410614
rect 591422 410378 591658 410614
rect 591102 410058 591338 410294
rect 591422 410058 591658 410294
rect 591102 374378 591338 374614
rect 591422 374378 591658 374614
rect 591102 374058 591338 374294
rect 591422 374058 591658 374294
rect 591102 338378 591338 338614
rect 591422 338378 591658 338614
rect 591102 338058 591338 338294
rect 591422 338058 591658 338294
rect 591102 302378 591338 302614
rect 591422 302378 591658 302614
rect 591102 302058 591338 302294
rect 591422 302058 591658 302294
rect 591102 266378 591338 266614
rect 591422 266378 591658 266614
rect 591102 266058 591338 266294
rect 591422 266058 591658 266294
rect 591102 230378 591338 230614
rect 591422 230378 591658 230614
rect 591102 230058 591338 230294
rect 591422 230058 591658 230294
rect 591102 194378 591338 194614
rect 591422 194378 591658 194614
rect 591102 194058 591338 194294
rect 591422 194058 591658 194294
rect 591102 158378 591338 158614
rect 591422 158378 591658 158614
rect 591102 158058 591338 158294
rect 591422 158058 591658 158294
rect 591102 122378 591338 122614
rect 591422 122378 591658 122614
rect 591102 122058 591338 122294
rect 591422 122058 591658 122294
rect 591102 86378 591338 86614
rect 591422 86378 591658 86614
rect 591102 86058 591338 86294
rect 591422 86058 591658 86294
rect 591102 50378 591338 50614
rect 591422 50378 591658 50614
rect 591102 50058 591338 50294
rect 591422 50058 591658 50294
rect 591102 14378 591338 14614
rect 591422 14378 591658 14614
rect 591102 14058 591338 14294
rect 591422 14058 591658 14294
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 680378 592298 680614
rect 592382 680378 592618 680614
rect 592062 680058 592298 680294
rect 592382 680058 592618 680294
rect 592062 644378 592298 644614
rect 592382 644378 592618 644614
rect 592062 644058 592298 644294
rect 592382 644058 592618 644294
rect 592062 608378 592298 608614
rect 592382 608378 592618 608614
rect 592062 608058 592298 608294
rect 592382 608058 592618 608294
rect 592062 572378 592298 572614
rect 592382 572378 592618 572614
rect 592062 572058 592298 572294
rect 592382 572058 592618 572294
rect 592062 536378 592298 536614
rect 592382 536378 592618 536614
rect 592062 536058 592298 536294
rect 592382 536058 592618 536294
rect 592062 500378 592298 500614
rect 592382 500378 592618 500614
rect 592062 500058 592298 500294
rect 592382 500058 592618 500294
rect 592062 464378 592298 464614
rect 592382 464378 592618 464614
rect 592062 464058 592298 464294
rect 592382 464058 592618 464294
rect 592062 428378 592298 428614
rect 592382 428378 592618 428614
rect 592062 428058 592298 428294
rect 592382 428058 592618 428294
rect 592062 392378 592298 392614
rect 592382 392378 592618 392614
rect 592062 392058 592298 392294
rect 592382 392058 592618 392294
rect 592062 356378 592298 356614
rect 592382 356378 592618 356614
rect 592062 356058 592298 356294
rect 592382 356058 592618 356294
rect 592062 320378 592298 320614
rect 592382 320378 592618 320614
rect 592062 320058 592298 320294
rect 592382 320058 592618 320294
rect 592062 284378 592298 284614
rect 592382 284378 592618 284614
rect 592062 284058 592298 284294
rect 592382 284058 592618 284294
rect 592062 248378 592298 248614
rect 592382 248378 592618 248614
rect 592062 248058 592298 248294
rect 592382 248058 592618 248294
rect 592062 212378 592298 212614
rect 592382 212378 592618 212614
rect 592062 212058 592298 212294
rect 592382 212058 592618 212294
rect 592062 176378 592298 176614
rect 592382 176378 592618 176614
rect 592062 176058 592298 176294
rect 592382 176058 592618 176294
rect 592062 140378 592298 140614
rect 592382 140378 592618 140614
rect 592062 140058 592298 140294
rect 592382 140058 592618 140294
rect 592062 104378 592298 104614
rect 592382 104378 592618 104614
rect 592062 104058 592298 104294
rect 592382 104058 592618 104294
rect 592062 68378 592298 68614
rect 592382 68378 592618 68614
rect 592062 68058 592298 68294
rect 592382 68058 592618 68294
rect 592062 32378 592298 32614
rect 592382 32378 592618 32614
rect 592062 32058 592298 32294
rect 592382 32058 592618 32294
rect 570986 -7302 571222 -7066
rect 571306 -7302 571542 -7066
rect 570986 -7622 571222 -7386
rect 571306 -7622 571542 -7386
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 592650 698294
rect -8726 698026 592650 698058
rect -6806 694894 590730 694926
rect -6806 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 590730 694894
rect -6806 694574 590730 694658
rect -6806 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 590730 694574
rect -6806 694306 590730 694338
rect -4886 691174 588810 691206
rect -4886 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 588810 691174
rect -4886 690854 588810 690938
rect -4886 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 588810 690854
rect -4886 690586 588810 690618
rect -2966 687454 586890 687486
rect -2966 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 586890 687454
rect -2966 687134 586890 687218
rect -2966 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 586890 687134
rect -2966 686866 586890 686898
rect -8726 680614 592650 680646
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect -8726 680294 592650 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect -8726 680026 592650 680058
rect -6806 676894 590730 676926
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect -6806 676574 590730 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect -6806 676306 590730 676338
rect -4886 673174 588810 673206
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect -4886 672854 588810 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect -4886 672586 588810 672618
rect -2966 669454 586890 669486
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect -2966 669134 586890 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect -2966 668866 586890 668898
rect -8726 662614 592650 662646
rect -8726 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 592650 662294
rect -8726 662026 592650 662058
rect -6806 658894 590730 658926
rect -6806 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 590730 658894
rect -6806 658574 590730 658658
rect -6806 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 590730 658574
rect -6806 658306 590730 658338
rect -4886 655174 588810 655206
rect -4886 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 588810 655174
rect -4886 654854 588810 654938
rect -4886 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 588810 654854
rect -4886 654586 588810 654618
rect -2966 651454 586890 651486
rect -2966 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 586890 651454
rect -2966 651134 586890 651218
rect -2966 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 586890 651134
rect -2966 650866 586890 650898
rect -8726 644614 592650 644646
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect -8726 644294 592650 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect -8726 644026 592650 644058
rect -6806 640894 590730 640926
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect -6806 640574 590730 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect -6806 640306 590730 640338
rect -4886 637174 588810 637206
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect -4886 636854 588810 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect -4886 636586 588810 636618
rect -2966 633454 586890 633486
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect -2966 633134 586890 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect -2966 632866 586890 632898
rect -8726 626614 592650 626646
rect -8726 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 592650 626294
rect -8726 626026 592650 626058
rect -6806 622894 590730 622926
rect -6806 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 590730 622894
rect -6806 622574 590730 622658
rect -6806 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 590730 622574
rect -6806 622306 590730 622338
rect -4886 619174 588810 619206
rect -4886 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 588810 619174
rect -4886 618854 588810 618938
rect -4886 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 588810 618854
rect -4886 618586 588810 618618
rect -2966 615454 586890 615486
rect -2966 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 586890 615454
rect -2966 615134 586890 615218
rect -2966 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 586890 615134
rect -2966 614866 586890 614898
rect -8726 608614 592650 608646
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect -8726 608294 592650 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect -8726 608026 592650 608058
rect -6806 604894 590730 604926
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect -6806 604574 590730 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect -6806 604306 590730 604338
rect -4886 601174 588810 601206
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect -4886 600854 588810 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect -4886 600586 588810 600618
rect -2966 597454 586890 597486
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect -2966 597134 586890 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect -2966 596866 586890 596898
rect -8726 590614 592650 590646
rect -8726 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 592650 590294
rect -8726 590026 592650 590058
rect -6806 586894 590730 586926
rect -6806 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 590730 586894
rect -6806 586574 590730 586658
rect -6806 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 590730 586574
rect -6806 586306 590730 586338
rect -4886 583174 588810 583206
rect -4886 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 77546 583174
rect 77782 582938 77866 583174
rect 78102 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 588810 583174
rect -4886 582854 588810 582938
rect -4886 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 77546 582854
rect 77782 582618 77866 582854
rect 78102 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 588810 582854
rect -4886 582586 588810 582618
rect -2966 579454 586890 579486
rect -2966 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 586890 579454
rect -2966 579134 586890 579218
rect -2966 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 586890 579134
rect -2966 578866 586890 578898
rect -8726 572614 592650 572646
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect -8726 572294 592650 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect -8726 572026 592650 572058
rect -6806 568894 590730 568926
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect -6806 568574 590730 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect -6806 568306 590730 568338
rect -4886 565174 588810 565206
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect -4886 564854 588810 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect -4886 564586 588810 564618
rect -2966 561454 586890 561486
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect -2966 561134 586890 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect -2966 560866 586890 560898
rect -8726 554614 592650 554646
rect -8726 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 84986 554614
rect 85222 554378 85306 554614
rect 85542 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 84986 554294
rect 85222 554058 85306 554294
rect 85542 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 592650 554294
rect -8726 554026 592650 554058
rect -6806 550894 590730 550926
rect -6806 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 81266 550894
rect 81502 550658 81586 550894
rect 81822 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 590730 550894
rect -6806 550574 590730 550658
rect -6806 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 81266 550574
rect 81502 550338 81586 550574
rect 81822 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 590730 550574
rect -6806 550306 590730 550338
rect -4886 547174 588810 547206
rect -4886 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 77546 547174
rect 77782 546938 77866 547174
rect 78102 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 588810 547174
rect -4886 546854 588810 546938
rect -4886 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 77546 546854
rect 77782 546618 77866 546854
rect 78102 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 588810 546854
rect -4886 546586 588810 546618
rect -2966 543454 586890 543486
rect -2966 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 586890 543454
rect -2966 543134 586890 543218
rect -2966 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 586890 543134
rect -2966 542866 586890 542898
rect -8726 536614 592650 536646
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 210986 536614
rect 211222 536378 211306 536614
rect 211542 536378 246986 536614
rect 247222 536378 247306 536614
rect 247542 536378 282986 536614
rect 283222 536378 283306 536614
rect 283542 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 354986 536614
rect 355222 536378 355306 536614
rect 355542 536378 390986 536614
rect 391222 536378 391306 536614
rect 391542 536378 426986 536614
rect 427222 536378 427306 536614
rect 427542 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect -8726 536294 592650 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 210986 536294
rect 211222 536058 211306 536294
rect 211542 536058 246986 536294
rect 247222 536058 247306 536294
rect 247542 536058 282986 536294
rect 283222 536058 283306 536294
rect 283542 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 354986 536294
rect 355222 536058 355306 536294
rect 355542 536058 390986 536294
rect 391222 536058 391306 536294
rect 391542 536058 426986 536294
rect 427222 536058 427306 536294
rect 427542 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect -8726 536026 592650 536058
rect -6806 532894 590730 532926
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 207266 532894
rect 207502 532658 207586 532894
rect 207822 532658 243266 532894
rect 243502 532658 243586 532894
rect 243822 532658 279266 532894
rect 279502 532658 279586 532894
rect 279822 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 351266 532894
rect 351502 532658 351586 532894
rect 351822 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 423266 532894
rect 423502 532658 423586 532894
rect 423822 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect -6806 532574 590730 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 207266 532574
rect 207502 532338 207586 532574
rect 207822 532338 243266 532574
rect 243502 532338 243586 532574
rect 243822 532338 279266 532574
rect 279502 532338 279586 532574
rect 279822 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 351266 532574
rect 351502 532338 351586 532574
rect 351822 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 423266 532574
rect 423502 532338 423586 532574
rect 423822 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect -6806 532306 590730 532338
rect -4886 529174 588810 529206
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 203546 529174
rect 203782 528938 203866 529174
rect 204102 528938 239546 529174
rect 239782 528938 239866 529174
rect 240102 528938 275546 529174
rect 275782 528938 275866 529174
rect 276102 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 347546 529174
rect 347782 528938 347866 529174
rect 348102 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect -4886 528854 588810 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 203546 528854
rect 203782 528618 203866 528854
rect 204102 528618 239546 528854
rect 239782 528618 239866 528854
rect 240102 528618 275546 528854
rect 275782 528618 275866 528854
rect 276102 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 347546 528854
rect 347782 528618 347866 528854
rect 348102 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect -4886 528586 588810 528618
rect -2966 525454 586890 525486
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect -2966 525134 586890 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect -2966 524866 586890 524898
rect -8726 518614 592650 518646
rect -8726 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 592650 518294
rect -8726 518026 592650 518058
rect -6806 514894 590730 514926
rect -6806 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 590730 514894
rect -6806 514574 590730 514658
rect -6806 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 590730 514574
rect -6806 514306 590730 514338
rect -4886 511174 588810 511206
rect -4886 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 588810 511174
rect -4886 510854 588810 510938
rect -4886 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 588810 510854
rect -4886 510586 588810 510618
rect -2966 507454 586890 507486
rect -2966 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 586890 507454
rect -2966 507134 586890 507218
rect -2966 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 586890 507134
rect -2966 506866 586890 506898
rect -8726 500614 592650 500646
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 174986 500614
rect 175222 500378 175306 500614
rect 175542 500378 210986 500614
rect 211222 500378 211306 500614
rect 211542 500378 246986 500614
rect 247222 500378 247306 500614
rect 247542 500378 282986 500614
rect 283222 500378 283306 500614
rect 283542 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect -8726 500294 592650 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 174986 500294
rect 175222 500058 175306 500294
rect 175542 500058 210986 500294
rect 211222 500058 211306 500294
rect 211542 500058 246986 500294
rect 247222 500058 247306 500294
rect 247542 500058 282986 500294
rect 283222 500058 283306 500294
rect 283542 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect -8726 500026 592650 500058
rect -6806 496894 590730 496926
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 171266 496894
rect 171502 496658 171586 496894
rect 171822 496658 207266 496894
rect 207502 496658 207586 496894
rect 207822 496658 243266 496894
rect 243502 496658 243586 496894
rect 243822 496658 279266 496894
rect 279502 496658 279586 496894
rect 279822 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect -6806 496574 590730 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 171266 496574
rect 171502 496338 171586 496574
rect 171822 496338 207266 496574
rect 207502 496338 207586 496574
rect 207822 496338 243266 496574
rect 243502 496338 243586 496574
rect 243822 496338 279266 496574
rect 279502 496338 279586 496574
rect 279822 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect -6806 496306 590730 496338
rect -4886 493174 588810 493206
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 167546 493174
rect 167782 492938 167866 493174
rect 168102 492938 203546 493174
rect 203782 492938 203866 493174
rect 204102 492938 239546 493174
rect 239782 492938 239866 493174
rect 240102 492938 275546 493174
rect 275782 492938 275866 493174
rect 276102 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect -4886 492854 588810 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 167546 492854
rect 167782 492618 167866 492854
rect 168102 492618 203546 492854
rect 203782 492618 203866 492854
rect 204102 492618 239546 492854
rect 239782 492618 239866 492854
rect 240102 492618 275546 492854
rect 275782 492618 275866 492854
rect 276102 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect -4886 492586 588810 492618
rect -2966 489454 586890 489486
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect -2966 489134 586890 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect -2966 488866 586890 488898
rect -8726 482614 592650 482646
rect -8726 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 592650 482294
rect -8726 482026 592650 482058
rect -6806 478894 590730 478926
rect -6806 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 590730 478894
rect -6806 478574 590730 478658
rect -6806 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 590730 478574
rect -6806 478306 590730 478338
rect -4886 475174 588810 475206
rect -4886 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 588810 475174
rect -4886 474854 588810 474938
rect -4886 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 588810 474854
rect -4886 474586 588810 474618
rect -2966 471454 586890 471486
rect -2966 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 244250 471454
rect 244486 471218 274970 471454
rect 275206 471218 305690 471454
rect 305926 471218 336410 471454
rect 336646 471218 367130 471454
rect 367366 471218 397850 471454
rect 398086 471218 428570 471454
rect 428806 471218 459290 471454
rect 459526 471218 490010 471454
rect 490246 471218 520730 471454
rect 520966 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 586890 471454
rect -2966 471134 586890 471218
rect -2966 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 244250 471134
rect 244486 470898 274970 471134
rect 275206 470898 305690 471134
rect 305926 470898 336410 471134
rect 336646 470898 367130 471134
rect 367366 470898 397850 471134
rect 398086 470898 428570 471134
rect 428806 470898 459290 471134
rect 459526 470898 490010 471134
rect 490246 470898 520730 471134
rect 520966 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 586890 471134
rect -2966 470866 586890 470898
rect -8726 464614 592650 464646
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect -8726 464294 592650 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect -8726 464026 592650 464058
rect -6806 460894 590730 460926
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect -6806 460574 590730 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect -6806 460306 590730 460338
rect -4886 457174 588810 457206
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect -4886 456854 588810 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect -4886 456586 588810 456618
rect -2966 453454 586890 453486
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 50328 453454
rect 50564 453218 186056 453454
rect 186292 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 259610 453454
rect 259846 453218 290330 453454
rect 290566 453218 321050 453454
rect 321286 453218 351770 453454
rect 352006 453218 382490 453454
rect 382726 453218 413210 453454
rect 413446 453218 443930 453454
rect 444166 453218 474650 453454
rect 474886 453218 505370 453454
rect 505606 453218 536090 453454
rect 536326 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect -2966 453134 586890 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 50328 453134
rect 50564 452898 186056 453134
rect 186292 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 259610 453134
rect 259846 452898 290330 453134
rect 290566 452898 321050 453134
rect 321286 452898 351770 453134
rect 352006 452898 382490 453134
rect 382726 452898 413210 453134
rect 413446 452898 443930 453134
rect 444166 452898 474650 453134
rect 474886 452898 505370 453134
rect 505606 452898 536090 453134
rect 536326 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect -2966 452866 586890 452898
rect -8726 446614 592650 446646
rect -8726 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 192986 446614
rect 193222 446378 193306 446614
rect 193542 446378 228986 446614
rect 229222 446378 229306 446614
rect 229542 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 192986 446294
rect 193222 446058 193306 446294
rect 193542 446058 228986 446294
rect 229222 446058 229306 446294
rect 229542 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 592650 446294
rect -8726 446026 592650 446058
rect -6806 442894 590730 442926
rect -6806 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 225266 442894
rect 225502 442658 225586 442894
rect 225822 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 590730 442894
rect -6806 442574 590730 442658
rect -6806 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 225266 442574
rect 225502 442338 225586 442574
rect 225822 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 590730 442574
rect -6806 442306 590730 442338
rect -4886 439174 588810 439206
rect -4886 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 221546 439174
rect 221782 438938 221866 439174
rect 222102 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 588810 439174
rect -4886 438854 588810 438938
rect -4886 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 221546 438854
rect 221782 438618 221866 438854
rect 222102 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 588810 438854
rect -4886 438586 588810 438618
rect -2966 435454 586890 435486
rect -2966 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 51008 435454
rect 51244 435218 185376 435454
rect 185612 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 244250 435454
rect 244486 435218 274970 435454
rect 275206 435218 305690 435454
rect 305926 435218 336410 435454
rect 336646 435218 367130 435454
rect 367366 435218 397850 435454
rect 398086 435218 428570 435454
rect 428806 435218 459290 435454
rect 459526 435218 490010 435454
rect 490246 435218 520730 435454
rect 520966 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 586890 435454
rect -2966 435134 586890 435218
rect -2966 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 51008 435134
rect 51244 434898 185376 435134
rect 185612 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 244250 435134
rect 244486 434898 274970 435134
rect 275206 434898 305690 435134
rect 305926 434898 336410 435134
rect 336646 434898 367130 435134
rect 367366 434898 397850 435134
rect 398086 434898 428570 435134
rect 428806 434898 459290 435134
rect 459526 434898 490010 435134
rect 490246 434898 520730 435134
rect 520966 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 586890 435134
rect -2966 434866 586890 434898
rect -8726 428614 592650 428646
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 210986 428614
rect 211222 428378 211306 428614
rect 211542 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect -8726 428294 592650 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 210986 428294
rect 211222 428058 211306 428294
rect 211542 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect -8726 428026 592650 428058
rect -6806 424894 590730 424926
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 207266 424894
rect 207502 424658 207586 424894
rect 207822 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect -6806 424574 590730 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 207266 424574
rect 207502 424338 207586 424574
rect 207822 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect -6806 424306 590730 424338
rect -4886 421174 588810 421206
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 203546 421174
rect 203782 420938 203866 421174
rect 204102 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect -4886 420854 588810 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 203546 420854
rect 203782 420618 203866 420854
rect 204102 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect -4886 420586 588810 420618
rect -2966 417454 586890 417486
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 50328 417454
rect 50564 417218 186056 417454
rect 186292 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 259610 417454
rect 259846 417218 290330 417454
rect 290566 417218 321050 417454
rect 321286 417218 351770 417454
rect 352006 417218 382490 417454
rect 382726 417218 413210 417454
rect 413446 417218 443930 417454
rect 444166 417218 474650 417454
rect 474886 417218 505370 417454
rect 505606 417218 536090 417454
rect 536326 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect -2966 417134 586890 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 50328 417134
rect 50564 416898 186056 417134
rect 186292 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 259610 417134
rect 259846 416898 290330 417134
rect 290566 416898 321050 417134
rect 321286 416898 351770 417134
rect 352006 416898 382490 417134
rect 382726 416898 413210 417134
rect 413446 416898 443930 417134
rect 444166 416898 474650 417134
rect 474886 416898 505370 417134
rect 505606 416898 536090 417134
rect 536326 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect -2966 416866 586890 416898
rect -8726 410614 592650 410646
rect -8726 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 192986 410614
rect 193222 410378 193306 410614
rect 193542 410378 228986 410614
rect 229222 410378 229306 410614
rect 229542 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 192986 410294
rect 193222 410058 193306 410294
rect 193542 410058 228986 410294
rect 229222 410058 229306 410294
rect 229542 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 592650 410294
rect -8726 410026 592650 410058
rect -6806 406894 590730 406926
rect -6806 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 189266 406894
rect 189502 406658 189586 406894
rect 189822 406658 225266 406894
rect 225502 406658 225586 406894
rect 225822 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 590730 406894
rect -6806 406574 590730 406658
rect -6806 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 189266 406574
rect 189502 406338 189586 406574
rect 189822 406338 225266 406574
rect 225502 406338 225586 406574
rect 225822 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 590730 406574
rect -6806 406306 590730 406338
rect -4886 403174 588810 403206
rect -4886 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 221546 403174
rect 221782 402938 221866 403174
rect 222102 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 588810 403174
rect -4886 402854 588810 402938
rect -4886 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 221546 402854
rect 221782 402618 221866 402854
rect 222102 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 588810 402854
rect -4886 402586 588810 402618
rect -2966 399454 586890 399486
rect -2966 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 51008 399454
rect 51244 399218 185376 399454
rect 185612 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 244250 399454
rect 244486 399218 274970 399454
rect 275206 399218 305690 399454
rect 305926 399218 336410 399454
rect 336646 399218 367130 399454
rect 367366 399218 397850 399454
rect 398086 399218 428570 399454
rect 428806 399218 459290 399454
rect 459526 399218 490010 399454
rect 490246 399218 520730 399454
rect 520966 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 586890 399454
rect -2966 399134 586890 399218
rect -2966 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 51008 399134
rect 51244 398898 185376 399134
rect 185612 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 244250 399134
rect 244486 398898 274970 399134
rect 275206 398898 305690 399134
rect 305926 398898 336410 399134
rect 336646 398898 367130 399134
rect 367366 398898 397850 399134
rect 398086 398898 428570 399134
rect 428806 398898 459290 399134
rect 459526 398898 490010 399134
rect 490246 398898 520730 399134
rect 520966 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 586890 399134
rect -2966 398866 586890 398898
rect -8726 392614 592650 392646
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 210986 392614
rect 211222 392378 211306 392614
rect 211542 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect -8726 392294 592650 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 210986 392294
rect 211222 392058 211306 392294
rect 211542 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect -8726 392026 592650 392058
rect -6806 388894 590730 388926
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 207266 388894
rect 207502 388658 207586 388894
rect 207822 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect -6806 388574 590730 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 207266 388574
rect 207502 388338 207586 388574
rect 207822 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect -6806 388306 590730 388338
rect -4886 385174 588810 385206
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 203546 385174
rect 203782 384938 203866 385174
rect 204102 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect -4886 384854 588810 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 203546 384854
rect 203782 384618 203866 384854
rect 204102 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect -4886 384586 588810 384618
rect -2966 381454 586890 381486
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 50328 381454
rect 50564 381218 186056 381454
rect 186292 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 259610 381454
rect 259846 381218 290330 381454
rect 290566 381218 321050 381454
rect 321286 381218 351770 381454
rect 352006 381218 382490 381454
rect 382726 381218 413210 381454
rect 413446 381218 443930 381454
rect 444166 381218 474650 381454
rect 474886 381218 505370 381454
rect 505606 381218 536090 381454
rect 536326 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect -2966 381134 586890 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 50328 381134
rect 50564 380898 186056 381134
rect 186292 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 259610 381134
rect 259846 380898 290330 381134
rect 290566 380898 321050 381134
rect 321286 380898 351770 381134
rect 352006 380898 382490 381134
rect 382726 380898 413210 381134
rect 413446 380898 443930 381134
rect 444166 380898 474650 381134
rect 474886 380898 505370 381134
rect 505606 380898 536090 381134
rect 536326 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect -2966 380866 586890 380898
rect -8726 374614 592650 374646
rect -8726 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 592650 374294
rect -8726 374026 592650 374058
rect -6806 370894 590730 370926
rect -6806 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 590730 370894
rect -6806 370574 590730 370658
rect -6806 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 590730 370574
rect -6806 370306 590730 370338
rect -4886 367174 588810 367206
rect -4886 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 588810 367174
rect -4886 366854 588810 366938
rect -4886 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 588810 366854
rect -4886 366586 588810 366618
rect -2966 363454 586890 363486
rect -2966 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 244250 363454
rect 244486 363218 274970 363454
rect 275206 363218 305690 363454
rect 305926 363218 336410 363454
rect 336646 363218 367130 363454
rect 367366 363218 397850 363454
rect 398086 363218 428570 363454
rect 428806 363218 459290 363454
rect 459526 363218 490010 363454
rect 490246 363218 520730 363454
rect 520966 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 586890 363454
rect -2966 363134 586890 363218
rect -2966 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 244250 363134
rect 244486 362898 274970 363134
rect 275206 362898 305690 363134
rect 305926 362898 336410 363134
rect 336646 362898 367130 363134
rect 367366 362898 397850 363134
rect 398086 362898 428570 363134
rect 428806 362898 459290 363134
rect 459526 362898 490010 363134
rect 490246 362898 520730 363134
rect 520966 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 586890 363134
rect -2966 362866 586890 362898
rect -8726 356614 592650 356646
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 102986 356614
rect 103222 356378 103306 356614
rect 103542 356378 138986 356614
rect 139222 356378 139306 356614
rect 139542 356378 174986 356614
rect 175222 356378 175306 356614
rect 175542 356378 210986 356614
rect 211222 356378 211306 356614
rect 211542 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect -8726 356294 592650 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 102986 356294
rect 103222 356058 103306 356294
rect 103542 356058 138986 356294
rect 139222 356058 139306 356294
rect 139542 356058 174986 356294
rect 175222 356058 175306 356294
rect 175542 356058 210986 356294
rect 211222 356058 211306 356294
rect 211542 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect -8726 356026 592650 356058
rect -6806 352894 590730 352926
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 63266 352894
rect 63502 352658 63586 352894
rect 63822 352658 99266 352894
rect 99502 352658 99586 352894
rect 99822 352658 135266 352894
rect 135502 352658 135586 352894
rect 135822 352658 171266 352894
rect 171502 352658 171586 352894
rect 171822 352658 207266 352894
rect 207502 352658 207586 352894
rect 207822 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect -6806 352574 590730 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 63266 352574
rect 63502 352338 63586 352574
rect 63822 352338 99266 352574
rect 99502 352338 99586 352574
rect 99822 352338 135266 352574
rect 135502 352338 135586 352574
rect 135822 352338 171266 352574
rect 171502 352338 171586 352574
rect 171822 352338 207266 352574
rect 207502 352338 207586 352574
rect 207822 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect -6806 352306 590730 352338
rect -4886 349174 588810 349206
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 59546 349174
rect 59782 348938 59866 349174
rect 60102 348938 95546 349174
rect 95782 348938 95866 349174
rect 96102 348938 131546 349174
rect 131782 348938 131866 349174
rect 132102 348938 167546 349174
rect 167782 348938 167866 349174
rect 168102 348938 203546 349174
rect 203782 348938 203866 349174
rect 204102 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect -4886 348854 588810 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 59546 348854
rect 59782 348618 59866 348854
rect 60102 348618 95546 348854
rect 95782 348618 95866 348854
rect 96102 348618 131546 348854
rect 131782 348618 131866 348854
rect 132102 348618 167546 348854
rect 167782 348618 167866 348854
rect 168102 348618 203546 348854
rect 203782 348618 203866 348854
rect 204102 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect -4886 348586 588810 348618
rect -2966 345454 586890 345486
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 259610 345454
rect 259846 345218 290330 345454
rect 290566 345218 321050 345454
rect 321286 345218 351770 345454
rect 352006 345218 382490 345454
rect 382726 345218 413210 345454
rect 413446 345218 443930 345454
rect 444166 345218 474650 345454
rect 474886 345218 505370 345454
rect 505606 345218 536090 345454
rect 536326 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect -2966 345134 586890 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 259610 345134
rect 259846 344898 290330 345134
rect 290566 344898 321050 345134
rect 321286 344898 351770 345134
rect 352006 344898 382490 345134
rect 382726 344898 413210 345134
rect 413446 344898 443930 345134
rect 444166 344898 474650 345134
rect 474886 344898 505370 345134
rect 505606 344898 536090 345134
rect 536326 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect -2966 344866 586890 344898
rect -8726 338614 592650 338646
rect -8726 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 84986 338614
rect 85222 338378 85306 338614
rect 85542 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 192986 338614
rect 193222 338378 193306 338614
rect 193542 338378 228986 338614
rect 229222 338378 229306 338614
rect 229542 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 84986 338294
rect 85222 338058 85306 338294
rect 85542 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 192986 338294
rect 193222 338058 193306 338294
rect 193542 338058 228986 338294
rect 229222 338058 229306 338294
rect 229542 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 592650 338294
rect -8726 338026 592650 338058
rect -6806 334894 590730 334926
rect -6806 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 189266 334894
rect 189502 334658 189586 334894
rect 189822 334658 225266 334894
rect 225502 334658 225586 334894
rect 225822 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 590730 334894
rect -6806 334574 590730 334658
rect -6806 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 189266 334574
rect 189502 334338 189586 334574
rect 189822 334338 225266 334574
rect 225502 334338 225586 334574
rect 225822 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 590730 334574
rect -6806 334306 590730 334338
rect -4886 331174 588810 331206
rect -4886 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 113546 331174
rect 113782 330938 113866 331174
rect 114102 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 221546 331174
rect 221782 330938 221866 331174
rect 222102 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 588810 331174
rect -4886 330854 588810 330938
rect -4886 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 113546 330854
rect 113782 330618 113866 330854
rect 114102 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 221546 330854
rect 221782 330618 221866 330854
rect 222102 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 588810 330854
rect -4886 330586 588810 330618
rect -2966 327454 586890 327486
rect -2966 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 244250 327454
rect 244486 327218 274970 327454
rect 275206 327218 305690 327454
rect 305926 327218 336410 327454
rect 336646 327218 367130 327454
rect 367366 327218 397850 327454
rect 398086 327218 428570 327454
rect 428806 327218 459290 327454
rect 459526 327218 490010 327454
rect 490246 327218 520730 327454
rect 520966 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 586890 327454
rect -2966 327134 586890 327218
rect -2966 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 244250 327134
rect 244486 326898 274970 327134
rect 275206 326898 305690 327134
rect 305926 326898 336410 327134
rect 336646 326898 367130 327134
rect 367366 326898 397850 327134
rect 398086 326898 428570 327134
rect 428806 326898 459290 327134
rect 459526 326898 490010 327134
rect 490246 326898 520730 327134
rect 520966 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 586890 327134
rect -2966 326866 586890 326898
rect -8726 320614 592650 320646
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 66986 320614
rect 67222 320378 67306 320614
rect 67542 320378 102986 320614
rect 103222 320378 103306 320614
rect 103542 320378 138986 320614
rect 139222 320378 139306 320614
rect 139542 320378 174986 320614
rect 175222 320378 175306 320614
rect 175542 320378 210986 320614
rect 211222 320378 211306 320614
rect 211542 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect -8726 320294 592650 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 66986 320294
rect 67222 320058 67306 320294
rect 67542 320058 102986 320294
rect 103222 320058 103306 320294
rect 103542 320058 138986 320294
rect 139222 320058 139306 320294
rect 139542 320058 174986 320294
rect 175222 320058 175306 320294
rect 175542 320058 210986 320294
rect 211222 320058 211306 320294
rect 211542 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect -8726 320026 592650 320058
rect -6806 316894 590730 316926
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 63266 316894
rect 63502 316658 63586 316894
rect 63822 316658 99266 316894
rect 99502 316658 99586 316894
rect 99822 316658 135266 316894
rect 135502 316658 135586 316894
rect 135822 316658 171266 316894
rect 171502 316658 171586 316894
rect 171822 316658 207266 316894
rect 207502 316658 207586 316894
rect 207822 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect -6806 316574 590730 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 63266 316574
rect 63502 316338 63586 316574
rect 63822 316338 99266 316574
rect 99502 316338 99586 316574
rect 99822 316338 135266 316574
rect 135502 316338 135586 316574
rect 135822 316338 171266 316574
rect 171502 316338 171586 316574
rect 171822 316338 207266 316574
rect 207502 316338 207586 316574
rect 207822 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect -6806 316306 590730 316338
rect -4886 313174 588810 313206
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 59546 313174
rect 59782 312938 59866 313174
rect 60102 312938 95546 313174
rect 95782 312938 95866 313174
rect 96102 312938 131546 313174
rect 131782 312938 131866 313174
rect 132102 312938 167546 313174
rect 167782 312938 167866 313174
rect 168102 312938 203546 313174
rect 203782 312938 203866 313174
rect 204102 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect -4886 312854 588810 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 59546 312854
rect 59782 312618 59866 312854
rect 60102 312618 95546 312854
rect 95782 312618 95866 312854
rect 96102 312618 131546 312854
rect 131782 312618 131866 312854
rect 132102 312618 167546 312854
rect 167782 312618 167866 312854
rect 168102 312618 203546 312854
rect 203782 312618 203866 312854
rect 204102 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect -4886 312586 588810 312618
rect -2966 309454 586890 309486
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 259610 309454
rect 259846 309218 290330 309454
rect 290566 309218 321050 309454
rect 321286 309218 351770 309454
rect 352006 309218 382490 309454
rect 382726 309218 413210 309454
rect 413446 309218 443930 309454
rect 444166 309218 474650 309454
rect 474886 309218 505370 309454
rect 505606 309218 536090 309454
rect 536326 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect -2966 309134 586890 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 259610 309134
rect 259846 308898 290330 309134
rect 290566 308898 321050 309134
rect 321286 308898 351770 309134
rect 352006 308898 382490 309134
rect 382726 308898 413210 309134
rect 413446 308898 443930 309134
rect 444166 308898 474650 309134
rect 474886 308898 505370 309134
rect 505606 308898 536090 309134
rect 536326 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect -2966 308866 586890 308898
rect -8726 302614 592650 302646
rect -8726 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 84986 302614
rect 85222 302378 85306 302614
rect 85542 302378 120986 302614
rect 121222 302378 121306 302614
rect 121542 302378 156986 302614
rect 157222 302378 157306 302614
rect 157542 302378 192986 302614
rect 193222 302378 193306 302614
rect 193542 302378 228986 302614
rect 229222 302378 229306 302614
rect 229542 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 84986 302294
rect 85222 302058 85306 302294
rect 85542 302058 120986 302294
rect 121222 302058 121306 302294
rect 121542 302058 156986 302294
rect 157222 302058 157306 302294
rect 157542 302058 192986 302294
rect 193222 302058 193306 302294
rect 193542 302058 228986 302294
rect 229222 302058 229306 302294
rect 229542 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 592650 302294
rect -8726 302026 592650 302058
rect -6806 298894 590730 298926
rect -6806 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 81266 298894
rect 81502 298658 81586 298894
rect 81822 298658 117266 298894
rect 117502 298658 117586 298894
rect 117822 298658 153266 298894
rect 153502 298658 153586 298894
rect 153822 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 225266 298894
rect 225502 298658 225586 298894
rect 225822 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 590730 298894
rect -6806 298574 590730 298658
rect -6806 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 81266 298574
rect 81502 298338 81586 298574
rect 81822 298338 117266 298574
rect 117502 298338 117586 298574
rect 117822 298338 153266 298574
rect 153502 298338 153586 298574
rect 153822 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 225266 298574
rect 225502 298338 225586 298574
rect 225822 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 590730 298574
rect -6806 298306 590730 298338
rect -4886 295174 588810 295206
rect -4886 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 77546 295174
rect 77782 294938 77866 295174
rect 78102 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 149546 295174
rect 149782 294938 149866 295174
rect 150102 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 221546 295174
rect 221782 294938 221866 295174
rect 222102 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 588810 295174
rect -4886 294854 588810 294938
rect -4886 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 77546 294854
rect 77782 294618 77866 294854
rect 78102 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 149546 294854
rect 149782 294618 149866 294854
rect 150102 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 221546 294854
rect 221782 294618 221866 294854
rect 222102 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 588810 294854
rect -4886 294586 588810 294618
rect -2966 291454 586890 291486
rect -2966 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 244250 291454
rect 244486 291218 274970 291454
rect 275206 291218 305690 291454
rect 305926 291218 336410 291454
rect 336646 291218 367130 291454
rect 367366 291218 397850 291454
rect 398086 291218 428570 291454
rect 428806 291218 459290 291454
rect 459526 291218 490010 291454
rect 490246 291218 520730 291454
rect 520966 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 586890 291454
rect -2966 291134 586890 291218
rect -2966 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 244250 291134
rect 244486 290898 274970 291134
rect 275206 290898 305690 291134
rect 305926 290898 336410 291134
rect 336646 290898 367130 291134
rect 367366 290898 397850 291134
rect 398086 290898 428570 291134
rect 428806 290898 459290 291134
rect 459526 290898 490010 291134
rect 490246 290898 520730 291134
rect 520966 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 586890 291134
rect -2966 290866 586890 290898
rect -8726 284614 592650 284646
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 210986 284614
rect 211222 284378 211306 284614
rect 211542 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect -8726 284294 592650 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 210986 284294
rect 211222 284058 211306 284294
rect 211542 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect -8726 284026 592650 284058
rect -6806 280894 590730 280926
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 207266 280894
rect 207502 280658 207586 280894
rect 207822 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect -6806 280574 590730 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 207266 280574
rect 207502 280338 207586 280574
rect 207822 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect -6806 280306 590730 280338
rect -4886 277174 588810 277206
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 203546 277174
rect 203782 276938 203866 277174
rect 204102 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect -4886 276854 588810 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 203546 276854
rect 203782 276618 203866 276854
rect 204102 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect -4886 276586 588810 276618
rect -2966 273454 586890 273486
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 50328 273454
rect 50564 273218 186056 273454
rect 186292 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 259610 273454
rect 259846 273218 290330 273454
rect 290566 273218 321050 273454
rect 321286 273218 351770 273454
rect 352006 273218 382490 273454
rect 382726 273218 413210 273454
rect 413446 273218 443930 273454
rect 444166 273218 474650 273454
rect 474886 273218 505370 273454
rect 505606 273218 536090 273454
rect 536326 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect -2966 273134 586890 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 50328 273134
rect 50564 272898 186056 273134
rect 186292 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 259610 273134
rect 259846 272898 290330 273134
rect 290566 272898 321050 273134
rect 321286 272898 351770 273134
rect 352006 272898 382490 273134
rect 382726 272898 413210 273134
rect 413446 272898 443930 273134
rect 444166 272898 474650 273134
rect 474886 272898 505370 273134
rect 505606 272898 536090 273134
rect 536326 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect -2966 272866 586890 272898
rect -8726 266614 592650 266646
rect -8726 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 192986 266614
rect 193222 266378 193306 266614
rect 193542 266378 228986 266614
rect 229222 266378 229306 266614
rect 229542 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 192986 266294
rect 193222 266058 193306 266294
rect 193542 266058 228986 266294
rect 229222 266058 229306 266294
rect 229542 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 592650 266294
rect -8726 266026 592650 266058
rect -6806 262894 590730 262926
rect -6806 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 225266 262894
rect 225502 262658 225586 262894
rect 225822 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 590730 262894
rect -6806 262574 590730 262658
rect -6806 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 225266 262574
rect 225502 262338 225586 262574
rect 225822 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 590730 262574
rect -6806 262306 590730 262338
rect -4886 259174 588810 259206
rect -4886 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 221546 259174
rect 221782 258938 221866 259174
rect 222102 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 588810 259174
rect -4886 258854 588810 258938
rect -4886 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 221546 258854
rect 221782 258618 221866 258854
rect 222102 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 588810 258854
rect -4886 258586 588810 258618
rect -2966 255454 586890 255486
rect -2966 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 51008 255454
rect 51244 255218 185376 255454
rect 185612 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 244250 255454
rect 244486 255218 274970 255454
rect 275206 255218 305690 255454
rect 305926 255218 336410 255454
rect 336646 255218 367130 255454
rect 367366 255218 397850 255454
rect 398086 255218 428570 255454
rect 428806 255218 459290 255454
rect 459526 255218 490010 255454
rect 490246 255218 520730 255454
rect 520966 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 586890 255454
rect -2966 255134 586890 255218
rect -2966 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 51008 255134
rect 51244 254898 185376 255134
rect 185612 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 244250 255134
rect 244486 254898 274970 255134
rect 275206 254898 305690 255134
rect 305926 254898 336410 255134
rect 336646 254898 367130 255134
rect 367366 254898 397850 255134
rect 398086 254898 428570 255134
rect 428806 254898 459290 255134
rect 459526 254898 490010 255134
rect 490246 254898 520730 255134
rect 520966 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 586890 255134
rect -2966 254866 586890 254898
rect -8726 248614 592650 248646
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 210986 248614
rect 211222 248378 211306 248614
rect 211542 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect -8726 248294 592650 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 210986 248294
rect 211222 248058 211306 248294
rect 211542 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect -8726 248026 592650 248058
rect -6806 244894 590730 244926
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 207266 244894
rect 207502 244658 207586 244894
rect 207822 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect -6806 244574 590730 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 207266 244574
rect 207502 244338 207586 244574
rect 207822 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect -6806 244306 590730 244338
rect -4886 241174 588810 241206
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 203546 241174
rect 203782 240938 203866 241174
rect 204102 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect -4886 240854 588810 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 203546 240854
rect 203782 240618 203866 240854
rect 204102 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect -4886 240586 588810 240618
rect -2966 237454 586890 237486
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 50328 237454
rect 50564 237218 186056 237454
rect 186292 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 259610 237454
rect 259846 237218 290330 237454
rect 290566 237218 321050 237454
rect 321286 237218 351770 237454
rect 352006 237218 382490 237454
rect 382726 237218 413210 237454
rect 413446 237218 443930 237454
rect 444166 237218 474650 237454
rect 474886 237218 505370 237454
rect 505606 237218 536090 237454
rect 536326 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect -2966 237134 586890 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 50328 237134
rect 50564 236898 186056 237134
rect 186292 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 259610 237134
rect 259846 236898 290330 237134
rect 290566 236898 321050 237134
rect 321286 236898 351770 237134
rect 352006 236898 382490 237134
rect 382726 236898 413210 237134
rect 413446 236898 443930 237134
rect 444166 236898 474650 237134
rect 474886 236898 505370 237134
rect 505606 236898 536090 237134
rect 536326 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect -2966 236866 586890 236898
rect -8726 230614 592650 230646
rect -8726 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 192986 230614
rect 193222 230378 193306 230614
rect 193542 230378 228986 230614
rect 229222 230378 229306 230614
rect 229542 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 192986 230294
rect 193222 230058 193306 230294
rect 193542 230058 228986 230294
rect 229222 230058 229306 230294
rect 229542 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 592650 230294
rect -8726 230026 592650 230058
rect -6806 226894 590730 226926
rect -6806 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 189266 226894
rect 189502 226658 189586 226894
rect 189822 226658 225266 226894
rect 225502 226658 225586 226894
rect 225822 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 590730 226894
rect -6806 226574 590730 226658
rect -6806 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 189266 226574
rect 189502 226338 189586 226574
rect 189822 226338 225266 226574
rect 225502 226338 225586 226574
rect 225822 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 590730 226574
rect -6806 226306 590730 226338
rect -4886 223174 588810 223206
rect -4886 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 221546 223174
rect 221782 222938 221866 223174
rect 222102 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 588810 223174
rect -4886 222854 588810 222938
rect -4886 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 221546 222854
rect 221782 222618 221866 222854
rect 222102 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 588810 222854
rect -4886 222586 588810 222618
rect -2966 219454 586890 219486
rect -2966 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 51008 219454
rect 51244 219218 185376 219454
rect 185612 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 244250 219454
rect 244486 219218 274970 219454
rect 275206 219218 305690 219454
rect 305926 219218 336410 219454
rect 336646 219218 367130 219454
rect 367366 219218 397850 219454
rect 398086 219218 428570 219454
rect 428806 219218 459290 219454
rect 459526 219218 490010 219454
rect 490246 219218 520730 219454
rect 520966 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 586890 219454
rect -2966 219134 586890 219218
rect -2966 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 51008 219134
rect 51244 218898 185376 219134
rect 185612 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 244250 219134
rect 244486 218898 274970 219134
rect 275206 218898 305690 219134
rect 305926 218898 336410 219134
rect 336646 218898 367130 219134
rect 367366 218898 397850 219134
rect 398086 218898 428570 219134
rect 428806 218898 459290 219134
rect 459526 218898 490010 219134
rect 490246 218898 520730 219134
rect 520966 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 586890 219134
rect -2966 218866 586890 218898
rect -8726 212614 592650 212646
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 210986 212614
rect 211222 212378 211306 212614
rect 211542 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect -8726 212294 592650 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 210986 212294
rect 211222 212058 211306 212294
rect 211542 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect -8726 212026 592650 212058
rect -6806 208894 590730 208926
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 207266 208894
rect 207502 208658 207586 208894
rect 207822 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect -6806 208574 590730 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 207266 208574
rect 207502 208338 207586 208574
rect 207822 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect -6806 208306 590730 208338
rect -4886 205174 588810 205206
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 203546 205174
rect 203782 204938 203866 205174
rect 204102 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect -4886 204854 588810 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 203546 204854
rect 203782 204618 203866 204854
rect 204102 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect -4886 204586 588810 204618
rect -2966 201454 586890 201486
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 50328 201454
rect 50564 201218 186056 201454
rect 186292 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 259610 201454
rect 259846 201218 290330 201454
rect 290566 201218 321050 201454
rect 321286 201218 351770 201454
rect 352006 201218 382490 201454
rect 382726 201218 413210 201454
rect 413446 201218 443930 201454
rect 444166 201218 474650 201454
rect 474886 201218 505370 201454
rect 505606 201218 536090 201454
rect 536326 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect -2966 201134 586890 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 50328 201134
rect 50564 200898 186056 201134
rect 186292 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 259610 201134
rect 259846 200898 290330 201134
rect 290566 200898 321050 201134
rect 321286 200898 351770 201134
rect 352006 200898 382490 201134
rect 382726 200898 413210 201134
rect 413446 200898 443930 201134
rect 444166 200898 474650 201134
rect 474886 200898 505370 201134
rect 505606 200898 536090 201134
rect 536326 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect -2966 200866 586890 200898
rect -8726 194614 592650 194646
rect -8726 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 120986 194614
rect 121222 194378 121306 194614
rect 121542 194378 156986 194614
rect 157222 194378 157306 194614
rect 157542 194378 192986 194614
rect 193222 194378 193306 194614
rect 193542 194378 228986 194614
rect 229222 194378 229306 194614
rect 229542 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 120986 194294
rect 121222 194058 121306 194294
rect 121542 194058 156986 194294
rect 157222 194058 157306 194294
rect 157542 194058 192986 194294
rect 193222 194058 193306 194294
rect 193542 194058 228986 194294
rect 229222 194058 229306 194294
rect 229542 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 592650 194294
rect -8726 194026 592650 194058
rect -6806 190894 590730 190926
rect -6806 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 117266 190894
rect 117502 190658 117586 190894
rect 117822 190658 153266 190894
rect 153502 190658 153586 190894
rect 153822 190658 189266 190894
rect 189502 190658 189586 190894
rect 189822 190658 225266 190894
rect 225502 190658 225586 190894
rect 225822 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 590730 190894
rect -6806 190574 590730 190658
rect -6806 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 117266 190574
rect 117502 190338 117586 190574
rect 117822 190338 153266 190574
rect 153502 190338 153586 190574
rect 153822 190338 189266 190574
rect 189502 190338 189586 190574
rect 189822 190338 225266 190574
rect 225502 190338 225586 190574
rect 225822 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 590730 190574
rect -6806 190306 590730 190338
rect -4886 187174 588810 187206
rect -4886 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 149546 187174
rect 149782 186938 149866 187174
rect 150102 186938 185546 187174
rect 185782 186938 185866 187174
rect 186102 186938 221546 187174
rect 221782 186938 221866 187174
rect 222102 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 588810 187174
rect -4886 186854 588810 186938
rect -4886 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 149546 186854
rect 149782 186618 149866 186854
rect 150102 186618 185546 186854
rect 185782 186618 185866 186854
rect 186102 186618 221546 186854
rect 221782 186618 221866 186854
rect 222102 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 588810 186854
rect -4886 186586 588810 186618
rect -2966 183454 586890 183486
rect -2966 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 244250 183454
rect 244486 183218 274970 183454
rect 275206 183218 305690 183454
rect 305926 183218 336410 183454
rect 336646 183218 367130 183454
rect 367366 183218 397850 183454
rect 398086 183218 428570 183454
rect 428806 183218 459290 183454
rect 459526 183218 490010 183454
rect 490246 183218 520730 183454
rect 520966 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 586890 183454
rect -2966 183134 586890 183218
rect -2966 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 244250 183134
rect 244486 182898 274970 183134
rect 275206 182898 305690 183134
rect 305926 182898 336410 183134
rect 336646 182898 367130 183134
rect 367366 182898 397850 183134
rect 398086 182898 428570 183134
rect 428806 182898 459290 183134
rect 459526 182898 490010 183134
rect 490246 182898 520730 183134
rect 520966 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 586890 183134
rect -2966 182866 586890 182898
rect -8726 176614 592650 176646
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 66986 176614
rect 67222 176378 67306 176614
rect 67542 176378 102986 176614
rect 103222 176378 103306 176614
rect 103542 176378 138986 176614
rect 139222 176378 139306 176614
rect 139542 176378 174986 176614
rect 175222 176378 175306 176614
rect 175542 176378 210986 176614
rect 211222 176378 211306 176614
rect 211542 176378 246986 176614
rect 247222 176378 247306 176614
rect 247542 176378 282986 176614
rect 283222 176378 283306 176614
rect 283542 176378 318986 176614
rect 319222 176378 319306 176614
rect 319542 176378 354986 176614
rect 355222 176378 355306 176614
rect 355542 176378 390986 176614
rect 391222 176378 391306 176614
rect 391542 176378 426986 176614
rect 427222 176378 427306 176614
rect 427542 176378 462986 176614
rect 463222 176378 463306 176614
rect 463542 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect -8726 176294 592650 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 66986 176294
rect 67222 176058 67306 176294
rect 67542 176058 102986 176294
rect 103222 176058 103306 176294
rect 103542 176058 138986 176294
rect 139222 176058 139306 176294
rect 139542 176058 174986 176294
rect 175222 176058 175306 176294
rect 175542 176058 210986 176294
rect 211222 176058 211306 176294
rect 211542 176058 246986 176294
rect 247222 176058 247306 176294
rect 247542 176058 282986 176294
rect 283222 176058 283306 176294
rect 283542 176058 318986 176294
rect 319222 176058 319306 176294
rect 319542 176058 354986 176294
rect 355222 176058 355306 176294
rect 355542 176058 390986 176294
rect 391222 176058 391306 176294
rect 391542 176058 426986 176294
rect 427222 176058 427306 176294
rect 427542 176058 462986 176294
rect 463222 176058 463306 176294
rect 463542 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect -8726 176026 592650 176058
rect -6806 172894 590730 172926
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 63266 172894
rect 63502 172658 63586 172894
rect 63822 172658 99266 172894
rect 99502 172658 99586 172894
rect 99822 172658 135266 172894
rect 135502 172658 135586 172894
rect 135822 172658 171266 172894
rect 171502 172658 171586 172894
rect 171822 172658 207266 172894
rect 207502 172658 207586 172894
rect 207822 172658 243266 172894
rect 243502 172658 243586 172894
rect 243822 172658 279266 172894
rect 279502 172658 279586 172894
rect 279822 172658 315266 172894
rect 315502 172658 315586 172894
rect 315822 172658 351266 172894
rect 351502 172658 351586 172894
rect 351822 172658 387266 172894
rect 387502 172658 387586 172894
rect 387822 172658 423266 172894
rect 423502 172658 423586 172894
rect 423822 172658 459266 172894
rect 459502 172658 459586 172894
rect 459822 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect -6806 172574 590730 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 63266 172574
rect 63502 172338 63586 172574
rect 63822 172338 99266 172574
rect 99502 172338 99586 172574
rect 99822 172338 135266 172574
rect 135502 172338 135586 172574
rect 135822 172338 171266 172574
rect 171502 172338 171586 172574
rect 171822 172338 207266 172574
rect 207502 172338 207586 172574
rect 207822 172338 243266 172574
rect 243502 172338 243586 172574
rect 243822 172338 279266 172574
rect 279502 172338 279586 172574
rect 279822 172338 315266 172574
rect 315502 172338 315586 172574
rect 315822 172338 351266 172574
rect 351502 172338 351586 172574
rect 351822 172338 387266 172574
rect 387502 172338 387586 172574
rect 387822 172338 423266 172574
rect 423502 172338 423586 172574
rect 423822 172338 459266 172574
rect 459502 172338 459586 172574
rect 459822 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect -6806 172306 590730 172338
rect -4886 169174 588810 169206
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 59546 169174
rect 59782 168938 59866 169174
rect 60102 168938 95546 169174
rect 95782 168938 95866 169174
rect 96102 168938 131546 169174
rect 131782 168938 131866 169174
rect 132102 168938 167546 169174
rect 167782 168938 167866 169174
rect 168102 168938 203546 169174
rect 203782 168938 203866 169174
rect 204102 168938 239546 169174
rect 239782 168938 239866 169174
rect 240102 168938 275546 169174
rect 275782 168938 275866 169174
rect 276102 168938 311546 169174
rect 311782 168938 311866 169174
rect 312102 168938 347546 169174
rect 347782 168938 347866 169174
rect 348102 168938 383546 169174
rect 383782 168938 383866 169174
rect 384102 168938 419546 169174
rect 419782 168938 419866 169174
rect 420102 168938 455546 169174
rect 455782 168938 455866 169174
rect 456102 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect -4886 168854 588810 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 59546 168854
rect 59782 168618 59866 168854
rect 60102 168618 95546 168854
rect 95782 168618 95866 168854
rect 96102 168618 131546 168854
rect 131782 168618 131866 168854
rect 132102 168618 167546 168854
rect 167782 168618 167866 168854
rect 168102 168618 203546 168854
rect 203782 168618 203866 168854
rect 204102 168618 239546 168854
rect 239782 168618 239866 168854
rect 240102 168618 275546 168854
rect 275782 168618 275866 168854
rect 276102 168618 311546 168854
rect 311782 168618 311866 168854
rect 312102 168618 347546 168854
rect 347782 168618 347866 168854
rect 348102 168618 383546 168854
rect 383782 168618 383866 168854
rect 384102 168618 419546 168854
rect 419782 168618 419866 168854
rect 420102 168618 455546 168854
rect 455782 168618 455866 168854
rect 456102 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect -4886 168586 588810 168618
rect -2966 165454 586890 165486
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 163826 165454
rect 164062 165218 164146 165454
rect 164382 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect -2966 165134 586890 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 163826 165134
rect 164062 164898 164146 165134
rect 164382 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect -2966 164866 586890 164898
rect -8726 158614 592650 158646
rect -8726 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 84986 158614
rect 85222 158378 85306 158614
rect 85542 158378 120986 158614
rect 121222 158378 121306 158614
rect 121542 158378 156986 158614
rect 157222 158378 157306 158614
rect 157542 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 228986 158614
rect 229222 158378 229306 158614
rect 229542 158378 264986 158614
rect 265222 158378 265306 158614
rect 265542 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 84986 158294
rect 85222 158058 85306 158294
rect 85542 158058 120986 158294
rect 121222 158058 121306 158294
rect 121542 158058 156986 158294
rect 157222 158058 157306 158294
rect 157542 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 228986 158294
rect 229222 158058 229306 158294
rect 229542 158058 264986 158294
rect 265222 158058 265306 158294
rect 265542 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 592650 158294
rect -8726 158026 592650 158058
rect -6806 154894 590730 154926
rect -6806 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 81266 154894
rect 81502 154658 81586 154894
rect 81822 154658 117266 154894
rect 117502 154658 117586 154894
rect 117822 154658 153266 154894
rect 153502 154658 153586 154894
rect 153822 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 225266 154894
rect 225502 154658 225586 154894
rect 225822 154658 261266 154894
rect 261502 154658 261586 154894
rect 261822 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 590730 154894
rect -6806 154574 590730 154658
rect -6806 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 81266 154574
rect 81502 154338 81586 154574
rect 81822 154338 117266 154574
rect 117502 154338 117586 154574
rect 117822 154338 153266 154574
rect 153502 154338 153586 154574
rect 153822 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 225266 154574
rect 225502 154338 225586 154574
rect 225822 154338 261266 154574
rect 261502 154338 261586 154574
rect 261822 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 590730 154574
rect -6806 154306 590730 154338
rect -4886 151174 588810 151206
rect -4886 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 77546 151174
rect 77782 150938 77866 151174
rect 78102 150938 113546 151174
rect 113782 150938 113866 151174
rect 114102 150938 149546 151174
rect 149782 150938 149866 151174
rect 150102 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 221546 151174
rect 221782 150938 221866 151174
rect 222102 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 588810 151174
rect -4886 150854 588810 150938
rect -4886 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 77546 150854
rect 77782 150618 77866 150854
rect 78102 150618 113546 150854
rect 113782 150618 113866 150854
rect 114102 150618 149546 150854
rect 149782 150618 149866 150854
rect 150102 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 221546 150854
rect 221782 150618 221866 150854
rect 222102 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 588810 150854
rect -4886 150586 588810 150618
rect -2966 147454 586890 147486
rect -2966 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 586890 147454
rect -2966 147134 586890 147218
rect -2966 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 586890 147134
rect -2966 146866 586890 146898
rect -8726 140614 592650 140646
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 66986 140614
rect 67222 140378 67306 140614
rect 67542 140378 102986 140614
rect 103222 140378 103306 140614
rect 103542 140378 138986 140614
rect 139222 140378 139306 140614
rect 139542 140378 174986 140614
rect 175222 140378 175306 140614
rect 175542 140378 210986 140614
rect 211222 140378 211306 140614
rect 211542 140378 246986 140614
rect 247222 140378 247306 140614
rect 247542 140378 282986 140614
rect 283222 140378 283306 140614
rect 283542 140378 318986 140614
rect 319222 140378 319306 140614
rect 319542 140378 354986 140614
rect 355222 140378 355306 140614
rect 355542 140378 390986 140614
rect 391222 140378 391306 140614
rect 391542 140378 426986 140614
rect 427222 140378 427306 140614
rect 427542 140378 462986 140614
rect 463222 140378 463306 140614
rect 463542 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect -8726 140294 592650 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 66986 140294
rect 67222 140058 67306 140294
rect 67542 140058 102986 140294
rect 103222 140058 103306 140294
rect 103542 140058 138986 140294
rect 139222 140058 139306 140294
rect 139542 140058 174986 140294
rect 175222 140058 175306 140294
rect 175542 140058 210986 140294
rect 211222 140058 211306 140294
rect 211542 140058 246986 140294
rect 247222 140058 247306 140294
rect 247542 140058 282986 140294
rect 283222 140058 283306 140294
rect 283542 140058 318986 140294
rect 319222 140058 319306 140294
rect 319542 140058 354986 140294
rect 355222 140058 355306 140294
rect 355542 140058 390986 140294
rect 391222 140058 391306 140294
rect 391542 140058 426986 140294
rect 427222 140058 427306 140294
rect 427542 140058 462986 140294
rect 463222 140058 463306 140294
rect 463542 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect -8726 140026 592650 140058
rect -6806 136894 590730 136926
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 99266 136894
rect 99502 136658 99586 136894
rect 99822 136658 135266 136894
rect 135502 136658 135586 136894
rect 135822 136658 171266 136894
rect 171502 136658 171586 136894
rect 171822 136658 207266 136894
rect 207502 136658 207586 136894
rect 207822 136658 243266 136894
rect 243502 136658 243586 136894
rect 243822 136658 279266 136894
rect 279502 136658 279586 136894
rect 279822 136658 315266 136894
rect 315502 136658 315586 136894
rect 315822 136658 351266 136894
rect 351502 136658 351586 136894
rect 351822 136658 387266 136894
rect 387502 136658 387586 136894
rect 387822 136658 423266 136894
rect 423502 136658 423586 136894
rect 423822 136658 459266 136894
rect 459502 136658 459586 136894
rect 459822 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect -6806 136574 590730 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 99266 136574
rect 99502 136338 99586 136574
rect 99822 136338 135266 136574
rect 135502 136338 135586 136574
rect 135822 136338 171266 136574
rect 171502 136338 171586 136574
rect 171822 136338 207266 136574
rect 207502 136338 207586 136574
rect 207822 136338 243266 136574
rect 243502 136338 243586 136574
rect 243822 136338 279266 136574
rect 279502 136338 279586 136574
rect 279822 136338 315266 136574
rect 315502 136338 315586 136574
rect 315822 136338 351266 136574
rect 351502 136338 351586 136574
rect 351822 136338 387266 136574
rect 387502 136338 387586 136574
rect 387822 136338 423266 136574
rect 423502 136338 423586 136574
rect 423822 136338 459266 136574
rect 459502 136338 459586 136574
rect 459822 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect -6806 136306 590730 136338
rect -4886 133174 588810 133206
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 95546 133174
rect 95782 132938 95866 133174
rect 96102 132938 131546 133174
rect 131782 132938 131866 133174
rect 132102 132938 167546 133174
rect 167782 132938 167866 133174
rect 168102 132938 203546 133174
rect 203782 132938 203866 133174
rect 204102 132938 239546 133174
rect 239782 132938 239866 133174
rect 240102 132938 275546 133174
rect 275782 132938 275866 133174
rect 276102 132938 311546 133174
rect 311782 132938 311866 133174
rect 312102 132938 347546 133174
rect 347782 132938 347866 133174
rect 348102 132938 383546 133174
rect 383782 132938 383866 133174
rect 384102 132938 419546 133174
rect 419782 132938 419866 133174
rect 420102 132938 455546 133174
rect 455782 132938 455866 133174
rect 456102 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect -4886 132854 588810 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 95546 132854
rect 95782 132618 95866 132854
rect 96102 132618 131546 132854
rect 131782 132618 131866 132854
rect 132102 132618 167546 132854
rect 167782 132618 167866 132854
rect 168102 132618 203546 132854
rect 203782 132618 203866 132854
rect 204102 132618 239546 132854
rect 239782 132618 239866 132854
rect 240102 132618 275546 132854
rect 275782 132618 275866 132854
rect 276102 132618 311546 132854
rect 311782 132618 311866 132854
rect 312102 132618 347546 132854
rect 347782 132618 347866 132854
rect 348102 132618 383546 132854
rect 383782 132618 383866 132854
rect 384102 132618 419546 132854
rect 419782 132618 419866 132854
rect 420102 132618 455546 132854
rect 455782 132618 455866 132854
rect 456102 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect -4886 132586 588810 132618
rect -2966 129454 586890 129486
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 127826 129454
rect 128062 129218 128146 129454
rect 128382 129218 163826 129454
rect 164062 129218 164146 129454
rect 164382 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect -2966 129134 586890 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 127826 129134
rect 128062 128898 128146 129134
rect 128382 128898 163826 129134
rect 164062 128898 164146 129134
rect 164382 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect -2966 128866 586890 128898
rect -8726 122614 592650 122646
rect -8726 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 84986 122614
rect 85222 122378 85306 122614
rect 85542 122378 120986 122614
rect 121222 122378 121306 122614
rect 121542 122378 156986 122614
rect 157222 122378 157306 122614
rect 157542 122378 192986 122614
rect 193222 122378 193306 122614
rect 193542 122378 228986 122614
rect 229222 122378 229306 122614
rect 229542 122378 264986 122614
rect 265222 122378 265306 122614
rect 265542 122378 300986 122614
rect 301222 122378 301306 122614
rect 301542 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 84986 122294
rect 85222 122058 85306 122294
rect 85542 122058 120986 122294
rect 121222 122058 121306 122294
rect 121542 122058 156986 122294
rect 157222 122058 157306 122294
rect 157542 122058 192986 122294
rect 193222 122058 193306 122294
rect 193542 122058 228986 122294
rect 229222 122058 229306 122294
rect 229542 122058 264986 122294
rect 265222 122058 265306 122294
rect 265542 122058 300986 122294
rect 301222 122058 301306 122294
rect 301542 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 592650 122294
rect -8726 122026 592650 122058
rect -6806 118894 590730 118926
rect -6806 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 81266 118894
rect 81502 118658 81586 118894
rect 81822 118658 117266 118894
rect 117502 118658 117586 118894
rect 117822 118658 153266 118894
rect 153502 118658 153586 118894
rect 153822 118658 189266 118894
rect 189502 118658 189586 118894
rect 189822 118658 225266 118894
rect 225502 118658 225586 118894
rect 225822 118658 261266 118894
rect 261502 118658 261586 118894
rect 261822 118658 297266 118894
rect 297502 118658 297586 118894
rect 297822 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 590730 118894
rect -6806 118574 590730 118658
rect -6806 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 81266 118574
rect 81502 118338 81586 118574
rect 81822 118338 117266 118574
rect 117502 118338 117586 118574
rect 117822 118338 153266 118574
rect 153502 118338 153586 118574
rect 153822 118338 189266 118574
rect 189502 118338 189586 118574
rect 189822 118338 225266 118574
rect 225502 118338 225586 118574
rect 225822 118338 261266 118574
rect 261502 118338 261586 118574
rect 261822 118338 297266 118574
rect 297502 118338 297586 118574
rect 297822 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 590730 118574
rect -6806 118306 590730 118338
rect -4886 115174 588810 115206
rect -4886 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 77546 115174
rect 77782 114938 77866 115174
rect 78102 114938 113546 115174
rect 113782 114938 113866 115174
rect 114102 114938 149546 115174
rect 149782 114938 149866 115174
rect 150102 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 221546 115174
rect 221782 114938 221866 115174
rect 222102 114938 257546 115174
rect 257782 114938 257866 115174
rect 258102 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 588810 115174
rect -4886 114854 588810 114938
rect -4886 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 77546 114854
rect 77782 114618 77866 114854
rect 78102 114618 113546 114854
rect 113782 114618 113866 114854
rect 114102 114618 149546 114854
rect 149782 114618 149866 114854
rect 150102 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 221546 114854
rect 221782 114618 221866 114854
rect 222102 114618 257546 114854
rect 257782 114618 257866 114854
rect 258102 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 588810 114854
rect -4886 114586 588810 114618
rect -2966 111454 586890 111486
rect -2966 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 586890 111454
rect -2966 111134 586890 111218
rect -2966 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 586890 111134
rect -2966 110866 586890 110898
rect -8726 104614 592650 104646
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 66986 104614
rect 67222 104378 67306 104614
rect 67542 104378 102986 104614
rect 103222 104378 103306 104614
rect 103542 104378 138986 104614
rect 139222 104378 139306 104614
rect 139542 104378 174986 104614
rect 175222 104378 175306 104614
rect 175542 104378 210986 104614
rect 211222 104378 211306 104614
rect 211542 104378 246986 104614
rect 247222 104378 247306 104614
rect 247542 104378 282986 104614
rect 283222 104378 283306 104614
rect 283542 104378 318986 104614
rect 319222 104378 319306 104614
rect 319542 104378 354986 104614
rect 355222 104378 355306 104614
rect 355542 104378 390986 104614
rect 391222 104378 391306 104614
rect 391542 104378 426986 104614
rect 427222 104378 427306 104614
rect 427542 104378 462986 104614
rect 463222 104378 463306 104614
rect 463542 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect -8726 104294 592650 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 66986 104294
rect 67222 104058 67306 104294
rect 67542 104058 102986 104294
rect 103222 104058 103306 104294
rect 103542 104058 138986 104294
rect 139222 104058 139306 104294
rect 139542 104058 174986 104294
rect 175222 104058 175306 104294
rect 175542 104058 210986 104294
rect 211222 104058 211306 104294
rect 211542 104058 246986 104294
rect 247222 104058 247306 104294
rect 247542 104058 282986 104294
rect 283222 104058 283306 104294
rect 283542 104058 318986 104294
rect 319222 104058 319306 104294
rect 319542 104058 354986 104294
rect 355222 104058 355306 104294
rect 355542 104058 390986 104294
rect 391222 104058 391306 104294
rect 391542 104058 426986 104294
rect 427222 104058 427306 104294
rect 427542 104058 462986 104294
rect 463222 104058 463306 104294
rect 463542 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect -8726 104026 592650 104058
rect -6806 100894 590730 100926
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 63266 100894
rect 63502 100658 63586 100894
rect 63822 100658 99266 100894
rect 99502 100658 99586 100894
rect 99822 100658 135266 100894
rect 135502 100658 135586 100894
rect 135822 100658 171266 100894
rect 171502 100658 171586 100894
rect 171822 100658 207266 100894
rect 207502 100658 207586 100894
rect 207822 100658 243266 100894
rect 243502 100658 243586 100894
rect 243822 100658 279266 100894
rect 279502 100658 279586 100894
rect 279822 100658 315266 100894
rect 315502 100658 315586 100894
rect 315822 100658 351266 100894
rect 351502 100658 351586 100894
rect 351822 100658 387266 100894
rect 387502 100658 387586 100894
rect 387822 100658 423266 100894
rect 423502 100658 423586 100894
rect 423822 100658 459266 100894
rect 459502 100658 459586 100894
rect 459822 100658 495266 100894
rect 495502 100658 495586 100894
rect 495822 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect -6806 100574 590730 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 63266 100574
rect 63502 100338 63586 100574
rect 63822 100338 99266 100574
rect 99502 100338 99586 100574
rect 99822 100338 135266 100574
rect 135502 100338 135586 100574
rect 135822 100338 171266 100574
rect 171502 100338 171586 100574
rect 171822 100338 207266 100574
rect 207502 100338 207586 100574
rect 207822 100338 243266 100574
rect 243502 100338 243586 100574
rect 243822 100338 279266 100574
rect 279502 100338 279586 100574
rect 279822 100338 315266 100574
rect 315502 100338 315586 100574
rect 315822 100338 351266 100574
rect 351502 100338 351586 100574
rect 351822 100338 387266 100574
rect 387502 100338 387586 100574
rect 387822 100338 423266 100574
rect 423502 100338 423586 100574
rect 423822 100338 459266 100574
rect 459502 100338 459586 100574
rect 459822 100338 495266 100574
rect 495502 100338 495586 100574
rect 495822 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect -6806 100306 590730 100338
rect -4886 97174 588810 97206
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 59546 97174
rect 59782 96938 59866 97174
rect 60102 96938 95546 97174
rect 95782 96938 95866 97174
rect 96102 96938 131546 97174
rect 131782 96938 131866 97174
rect 132102 96938 167546 97174
rect 167782 96938 167866 97174
rect 168102 96938 203546 97174
rect 203782 96938 203866 97174
rect 204102 96938 239546 97174
rect 239782 96938 239866 97174
rect 240102 96938 275546 97174
rect 275782 96938 275866 97174
rect 276102 96938 311546 97174
rect 311782 96938 311866 97174
rect 312102 96938 347546 97174
rect 347782 96938 347866 97174
rect 348102 96938 383546 97174
rect 383782 96938 383866 97174
rect 384102 96938 419546 97174
rect 419782 96938 419866 97174
rect 420102 96938 455546 97174
rect 455782 96938 455866 97174
rect 456102 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect -4886 96854 588810 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 59546 96854
rect 59782 96618 59866 96854
rect 60102 96618 95546 96854
rect 95782 96618 95866 96854
rect 96102 96618 131546 96854
rect 131782 96618 131866 96854
rect 132102 96618 167546 96854
rect 167782 96618 167866 96854
rect 168102 96618 203546 96854
rect 203782 96618 203866 96854
rect 204102 96618 239546 96854
rect 239782 96618 239866 96854
rect 240102 96618 275546 96854
rect 275782 96618 275866 96854
rect 276102 96618 311546 96854
rect 311782 96618 311866 96854
rect 312102 96618 347546 96854
rect 347782 96618 347866 96854
rect 348102 96618 383546 96854
rect 383782 96618 383866 96854
rect 384102 96618 419546 96854
rect 419782 96618 419866 96854
rect 420102 96618 455546 96854
rect 455782 96618 455866 96854
rect 456102 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect -4886 96586 588810 96618
rect -2966 93454 586890 93486
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 127826 93454
rect 128062 93218 128146 93454
rect 128382 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect -2966 93134 586890 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 127826 93134
rect 128062 92898 128146 93134
rect 128382 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect -2966 92866 586890 92898
rect -8726 86614 592650 86646
rect -8726 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 120986 86614
rect 121222 86378 121306 86614
rect 121542 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 192986 86614
rect 193222 86378 193306 86614
rect 193542 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 120986 86294
rect 121222 86058 121306 86294
rect 121542 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 192986 86294
rect 193222 86058 193306 86294
rect 193542 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 592650 86294
rect -8726 86026 592650 86058
rect -6806 82894 590730 82926
rect -6806 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 117266 82894
rect 117502 82658 117586 82894
rect 117822 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 189266 82894
rect 189502 82658 189586 82894
rect 189822 82658 225266 82894
rect 225502 82658 225586 82894
rect 225822 82658 261266 82894
rect 261502 82658 261586 82894
rect 261822 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 590730 82894
rect -6806 82574 590730 82658
rect -6806 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 117266 82574
rect 117502 82338 117586 82574
rect 117822 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 189266 82574
rect 189502 82338 189586 82574
rect 189822 82338 225266 82574
rect 225502 82338 225586 82574
rect 225822 82338 261266 82574
rect 261502 82338 261586 82574
rect 261822 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 590730 82574
rect -6806 82306 590730 82338
rect -4886 79174 588810 79206
rect -4886 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 588810 79174
rect -4886 78854 588810 78938
rect -4886 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 588810 78854
rect -4886 78586 588810 78618
rect -2966 75454 586890 75486
rect -2966 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 586890 75454
rect -2966 75134 586890 75218
rect -2966 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 586890 75134
rect -2966 74866 586890 74898
rect -8726 68614 592650 68646
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 66986 68614
rect 67222 68378 67306 68614
rect 67542 68378 102986 68614
rect 103222 68378 103306 68614
rect 103542 68378 138986 68614
rect 139222 68378 139306 68614
rect 139542 68378 174986 68614
rect 175222 68378 175306 68614
rect 175542 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 246986 68614
rect 247222 68378 247306 68614
rect 247542 68378 282986 68614
rect 283222 68378 283306 68614
rect 283542 68378 318986 68614
rect 319222 68378 319306 68614
rect 319542 68378 354986 68614
rect 355222 68378 355306 68614
rect 355542 68378 390986 68614
rect 391222 68378 391306 68614
rect 391542 68378 426986 68614
rect 427222 68378 427306 68614
rect 427542 68378 462986 68614
rect 463222 68378 463306 68614
rect 463542 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect -8726 68294 592650 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 66986 68294
rect 67222 68058 67306 68294
rect 67542 68058 102986 68294
rect 103222 68058 103306 68294
rect 103542 68058 138986 68294
rect 139222 68058 139306 68294
rect 139542 68058 174986 68294
rect 175222 68058 175306 68294
rect 175542 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 246986 68294
rect 247222 68058 247306 68294
rect 247542 68058 282986 68294
rect 283222 68058 283306 68294
rect 283542 68058 318986 68294
rect 319222 68058 319306 68294
rect 319542 68058 354986 68294
rect 355222 68058 355306 68294
rect 355542 68058 390986 68294
rect 391222 68058 391306 68294
rect 391542 68058 426986 68294
rect 427222 68058 427306 68294
rect 427542 68058 462986 68294
rect 463222 68058 463306 68294
rect 463542 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect -8726 68026 592650 68058
rect -6806 64894 590730 64926
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 63266 64894
rect 63502 64658 63586 64894
rect 63822 64658 99266 64894
rect 99502 64658 99586 64894
rect 99822 64658 135266 64894
rect 135502 64658 135586 64894
rect 135822 64658 171266 64894
rect 171502 64658 171586 64894
rect 171822 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 243266 64894
rect 243502 64658 243586 64894
rect 243822 64658 279266 64894
rect 279502 64658 279586 64894
rect 279822 64658 315266 64894
rect 315502 64658 315586 64894
rect 315822 64658 351266 64894
rect 351502 64658 351586 64894
rect 351822 64658 387266 64894
rect 387502 64658 387586 64894
rect 387822 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect -6806 64574 590730 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 63266 64574
rect 63502 64338 63586 64574
rect 63822 64338 99266 64574
rect 99502 64338 99586 64574
rect 99822 64338 135266 64574
rect 135502 64338 135586 64574
rect 135822 64338 171266 64574
rect 171502 64338 171586 64574
rect 171822 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 243266 64574
rect 243502 64338 243586 64574
rect 243822 64338 279266 64574
rect 279502 64338 279586 64574
rect 279822 64338 315266 64574
rect 315502 64338 315586 64574
rect 315822 64338 351266 64574
rect 351502 64338 351586 64574
rect 351822 64338 387266 64574
rect 387502 64338 387586 64574
rect 387822 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect -6806 64306 590730 64338
rect -4886 61174 588810 61206
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 59546 61174
rect 59782 60938 59866 61174
rect 60102 60938 95546 61174
rect 95782 60938 95866 61174
rect 96102 60938 131546 61174
rect 131782 60938 131866 61174
rect 132102 60938 167546 61174
rect 167782 60938 167866 61174
rect 168102 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 239546 61174
rect 239782 60938 239866 61174
rect 240102 60938 275546 61174
rect 275782 60938 275866 61174
rect 276102 60938 311546 61174
rect 311782 60938 311866 61174
rect 312102 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect -4886 60854 588810 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 59546 60854
rect 59782 60618 59866 60854
rect 60102 60618 95546 60854
rect 95782 60618 95866 60854
rect 96102 60618 131546 60854
rect 131782 60618 131866 60854
rect 132102 60618 167546 60854
rect 167782 60618 167866 60854
rect 168102 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 239546 60854
rect 239782 60618 239866 60854
rect 240102 60618 275546 60854
rect 275782 60618 275866 60854
rect 276102 60618 311546 60854
rect 311782 60618 311866 60854
rect 312102 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect -4886 60586 588810 60618
rect -2966 57454 586890 57486
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect -2966 57134 586890 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect -2966 56866 586890 56898
rect -8726 50614 592650 50646
rect -8726 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 592650 50294
rect -8726 50026 592650 50058
rect -6806 46894 590730 46926
rect -6806 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 590730 46894
rect -6806 46574 590730 46658
rect -6806 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 590730 46574
rect -6806 46306 590730 46338
rect -4886 43174 588810 43206
rect -4886 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 588810 43174
rect -4886 42854 588810 42938
rect -4886 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 588810 42854
rect -4886 42586 588810 42618
rect -2966 39454 586890 39486
rect -2966 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 586890 39454
rect -2966 39134 586890 39218
rect -2966 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 586890 39134
rect -2966 38866 586890 38898
rect -8726 32614 592650 32646
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect -8726 32294 592650 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect -8726 32026 592650 32058
rect -6806 28894 590730 28926
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect -6806 28574 590730 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect -6806 28306 590730 28338
rect -4886 25174 588810 25206
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect -4886 24854 588810 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect -4886 24586 588810 24618
rect -2966 21454 586890 21486
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect -2966 21134 586890 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect -2966 20866 586890 20898
rect -8726 14614 592650 14646
rect -8726 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 592650 14294
rect -8726 14026 592650 14058
rect -6806 10894 590730 10926
rect -6806 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 590730 10894
rect -6806 10574 590730 10658
rect -6806 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 590730 10574
rect -6806 10306 590730 10338
rect -4886 7174 588810 7206
rect -4886 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 588810 7174
rect -4886 6854 588810 6938
rect -4886 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 588810 6854
rect -4886 6586 588810 6618
rect -2966 3454 586890 3486
rect -2966 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 586890 3454
rect -2966 3134 586890 3218
rect -2966 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 586890 3134
rect -2966 2866 586890 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use sky130_sram_2kbyte_1rw1r_32x512_8  BB_SRAM
timestamp 0
transform 1 0 50000 0 1 380000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  VB_SRAM
timestamp 0
transform 1 0 50000 0 1 200000
box 0 0 136620 83308
use c0_system  mprj
timestamp 0
transform 1 0 240000 0 1 180000
box 0 0 298816 299464
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 38866 586890 39486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 74866 586890 75486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 110866 586890 111486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 146866 586890 147486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 182866 586890 183486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 218866 586890 219486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 254866 586890 255486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 290866 586890 291486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 326866 586890 327486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 362866 586890 363486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 398866 586890 399486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 434866 586890 435486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 470866 586890 471486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 578866 586890 579486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 614866 586890 615486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 650866 586890 651486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 686866 586890 687486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 -1894 254414 178000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 -1894 290414 178000 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 -1894 326414 178000 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 -1894 362414 178000 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 -1894 398414 178000 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 -1894 434414 178000 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 -1894 470414 178000 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 -1894 506414 178000 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 -1894 542414 178000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 -1894 74414 198000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 -1894 110414 198000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 -1894 146414 198000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 -1894 182414 198000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 285308 74414 378000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 285308 110414 378000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 285308 146414 378000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 285308 182414 378000 6 vccd1
port 531 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 1794 -1894 2414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 -1894 38414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 465308 74414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 465308 110414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 465308 146414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 465308 182414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 -1894 218414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 482000 254414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 482000 290414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 482000 326414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 482000 362414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 482000 398414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 482000 434414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 482000 470414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 482000 506414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 482000 542414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 577794 -1894 578414 705830 6 vccd1
port 531 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 532 nsew power input
rlabel metal5 s -4886 6586 588810 7206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 42586 588810 43206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 78586 588810 79206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 114586 588810 115206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 150586 588810 151206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 186586 588810 187206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 222586 588810 223206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 258586 588810 259206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 294586 588810 295206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 330586 588810 331206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 366586 588810 367206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 402586 588810 403206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 438586 588810 439206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 474586 588810 475206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 510586 588810 511206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 546586 588810 547206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 582586 588810 583206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 618586 588810 619206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 654586 588810 655206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 690586 588810 691206 6 vccd2
port 532 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 -3814 258134 178000 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 -3814 294134 178000 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 -3814 330134 178000 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 -3814 366134 178000 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 -3814 402134 178000 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 -3814 438134 178000 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 -3814 474134 178000 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 -3814 510134 178000 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 -3814 78134 198000 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 -3814 114134 198000 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 -3814 150134 198000 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 -3814 186134 198000 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 285308 78134 378000 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 285308 114134 378000 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 285308 150134 378000 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 285308 186134 378000 6 vccd2
port 532 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 532 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 5514 -3814 6134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 41514 -3814 42134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 465308 78134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 465308 114134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 465308 150134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 465308 186134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 -3814 222134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 482000 258134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 482000 294134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 482000 330134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 482000 366134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 482000 402134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 482000 438134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 482000 474134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 482000 510134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 545514 -3814 546134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 581514 -3814 582134 707750 6 vccd2
port 532 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 533 nsew power input
rlabel metal5 s -6806 10306 590730 10926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 46306 590730 46926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 82306 590730 82926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 118306 590730 118926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 154306 590730 154926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 190306 590730 190926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 226306 590730 226926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 262306 590730 262926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 298306 590730 298926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 334306 590730 334926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 370306 590730 370926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 406306 590730 406926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 442306 590730 442926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 478306 590730 478926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 514306 590730 514926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 550306 590730 550926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 586306 590730 586926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 622306 590730 622926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 658306 590730 658926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 694306 590730 694926 6 vdda1
port 533 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 -5734 261854 178000 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 -5734 297854 178000 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 -5734 333854 178000 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 -5734 369854 178000 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 -5734 405854 178000 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 -5734 441854 178000 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 -5734 477854 178000 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 -5734 513854 178000 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 -5734 81854 198000 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 -5734 117854 198000 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 -5734 153854 198000 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 285308 81854 378000 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 285308 117854 378000 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 285308 153854 378000 6 vdda1
port 533 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 533 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 9234 -5734 9854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 45234 -5734 45854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 465308 81854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 465308 117854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 465308 153854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 -5734 189854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 -5734 225854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 482000 261854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 482000 297854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 482000 333854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 482000 369854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 482000 405854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 482000 441854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 482000 477854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 482000 513854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 549234 -5734 549854 709670 6 vdda1
port 533 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 534 nsew power input
rlabel metal5 s -8726 14026 592650 14646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 50026 592650 50646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 86026 592650 86646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 122026 592650 122646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 158026 592650 158646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 194026 592650 194646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 230026 592650 230646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 266026 592650 266646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 302026 592650 302646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 338026 592650 338646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 374026 592650 374646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 410026 592650 410646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 446026 592650 446646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 482026 592650 482646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 518026 592650 518646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 554026 592650 554646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 590026 592650 590646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 626026 592650 626646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 662026 592650 662646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 698026 592650 698646 6 vdda2
port 534 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 -7654 265574 178000 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 -7654 301574 178000 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 -7654 337574 178000 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 -7654 373574 178000 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 -7654 409574 178000 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 -7654 445574 178000 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 -7654 481574 178000 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 -7654 517574 178000 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 -7654 49574 198000 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 -7654 85574 198000 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 -7654 121574 198000 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 -7654 157574 198000 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 285308 49574 378000 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 285308 85574 378000 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 285308 121574 378000 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 285308 157574 378000 6 vdda2
port 534 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 534 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 12954 -7654 13574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 465308 49574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 465308 85574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 465308 121574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 465308 157574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 -7654 193574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 -7654 229574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 482000 265574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 482000 301574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 482000 337574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 482000 373574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 482000 409574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 482000 445574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 482000 481574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 482000 517574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 552954 -7654 553574 711590 6 vdda2
port 534 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 28306 590730 28926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 64306 590730 64926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 100306 590730 100926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 136306 590730 136926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 172306 590730 172926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 208306 590730 208926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 244306 590730 244926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 280306 590730 280926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 316306 590730 316926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 352306 590730 352926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 388306 590730 388926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 424306 590730 424926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 460306 590730 460926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 496306 590730 496926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 532306 590730 532926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 568306 590730 568926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 604306 590730 604926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 640306 590730 640926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 676306 590730 676926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 -5734 243854 178000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 -5734 279854 178000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 -5734 315854 178000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 -5734 351854 178000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 -5734 387854 178000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 -5734 423854 178000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 -5734 459854 178000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 -5734 495854 178000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 -5734 531854 178000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 -5734 63854 198000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 -5734 99854 198000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 -5734 135854 198000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 -5734 171854 198000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 285308 63854 378000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 285308 99854 378000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 285308 135854 378000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 285308 171854 378000 6 vssa1
port 535 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 535 nsew ground input
rlabel metal4 s 27234 -5734 27854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 465308 63854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 465308 99854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 465308 135854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 465308 171854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 -5734 207854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 482000 243854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 482000 279854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 482000 315854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 482000 351854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 482000 387854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 482000 423854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 482000 459854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 482000 495854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 482000 531854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 567234 -5734 567854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 32026 592650 32646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 68026 592650 68646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 104026 592650 104646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 140026 592650 140646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 176026 592650 176646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 212026 592650 212646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 248026 592650 248646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 284026 592650 284646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 320026 592650 320646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 356026 592650 356646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 392026 592650 392646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 428026 592650 428646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 464026 592650 464646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 500026 592650 500646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 536026 592650 536646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 572026 592650 572646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 608026 592650 608646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 644026 592650 644646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 680026 592650 680646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 -7654 247574 178000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 -7654 283574 178000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 -7654 319574 178000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 -7654 355574 178000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 -7654 391574 178000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 -7654 427574 178000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 -7654 463574 178000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 -7654 499574 178000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 -7654 535574 178000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 -7654 67574 198000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 -7654 103574 198000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 -7654 139574 198000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 -7654 175574 198000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 285308 67574 378000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 285308 103574 378000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 285308 139574 378000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 285308 175574 378000 6 vssa2
port 536 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 -7654 31574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 465308 67574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 465308 103574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 465308 139574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 465308 175574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 -7654 211574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 482000 247574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 482000 283574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 482000 319574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 482000 355574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 482000 391574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 482000 427574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 482000 463574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 482000 499574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 482000 535574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 570954 -7654 571574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 20866 586890 21486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 56866 586890 57486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 92866 586890 93486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 128866 586890 129486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 164866 586890 165486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 200866 586890 201486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 236866 586890 237486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 272866 586890 273486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 308866 586890 309486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 344866 586890 345486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 380866 586890 381486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 416866 586890 417486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 452866 586890 453486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 488866 586890 489486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 524866 586890 525486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 560866 586890 561486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 596866 586890 597486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 632866 586890 633486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 668866 586890 669486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 -1894 272414 178000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 -1894 308414 178000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 -1894 344414 178000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 -1894 380414 178000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 -1894 416414 178000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 -1894 452414 178000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 -1894 488414 178000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 -1894 524414 178000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 -1894 56414 198000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 -1894 92414 198000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 -1894 128414 198000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 -1894 164414 198000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 285308 56414 378000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 285308 92414 378000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 285308 128414 378000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 285308 164414 378000 6 vssd1
port 537 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 537 nsew ground input
rlabel metal4 s 19794 -1894 20414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 465308 56414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 465308 92414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 465308 128414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 465308 164414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 -1894 200414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 -1894 236414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 482000 272414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 482000 308414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 482000 344414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 482000 380414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 482000 416414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 482000 452414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 482000 488414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 482000 524414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 559794 -1894 560414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 24586 588810 25206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 60586 588810 61206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 96586 588810 97206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 132586 588810 133206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 168586 588810 169206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 204586 588810 205206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 240586 588810 241206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 276586 588810 277206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 312586 588810 313206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 348586 588810 349206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 384586 588810 385206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 420586 588810 421206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 456586 588810 457206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 492586 588810 493206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 528586 588810 529206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 564586 588810 565206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 600586 588810 601206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 636586 588810 637206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 672586 588810 673206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 -3814 240134 178000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 -3814 276134 178000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 -3814 312134 178000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 -3814 348134 178000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 -3814 384134 178000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 -3814 420134 178000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 -3814 456134 178000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 -3814 492134 178000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 -3814 528134 178000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 -3814 60134 198000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 -3814 96134 198000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 -3814 132134 198000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 -3814 168134 198000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 285308 60134 378000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 285308 96134 378000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 285308 132134 378000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 285308 168134 378000 6 vssd2
port 538 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 538 nsew ground input
rlabel metal4 s 23514 -3814 24134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 465308 60134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 465308 96134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 465308 132134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 465308 168134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 -3814 204134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 482000 240134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 482000 276134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 482000 312134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 482000 348134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 482000 384134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 482000 420134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 482000 456134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 482000 492134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 482000 528134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 563514 -3814 564134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 541 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 607 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 608 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 609 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 610 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 611 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 612 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 613 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 614 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 615 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 616 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 617 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 618 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 619 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 620 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 621 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 622 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 623 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 624 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 625 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 626 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 627 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 628 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 629 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 630 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 631 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 632 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 633 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 634 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 635 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 636 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 637 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 638 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO c0_system
  CLASS BLOCK ;
  FOREIGN c0_system ;
  ORIGIN 0.000 0.000 ;
  SIZE 1200.000 BY 1800.000 ;
  PIN bb_addr0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 805.160 4.000 805.760 ;
    END
  END bb_addr0[0]
  PIN bb_addr0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1133.600 4.000 1134.200 ;
    END
  END bb_addr0[10]
  PIN bb_addr0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1164.200 4.000 1164.800 ;
    END
  END bb_addr0[11]
  PIN bb_addr0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1194.120 4.000 1194.720 ;
    END
  END bb_addr0[12]
  PIN bb_addr0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1224.720 4.000 1225.320 ;
    END
  END bb_addr0[13]
  PIN bb_addr0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1255.320 4.000 1255.920 ;
    END
  END bb_addr0[14]
  PIN bb_addr0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1285.240 4.000 1285.840 ;
    END
  END bb_addr0[15]
  PIN bb_addr0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1315.840 4.000 1316.440 ;
    END
  END bb_addr0[16]
  PIN bb_addr0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1346.440 4.000 1347.040 ;
    END
  END bb_addr0[17]
  PIN bb_addr0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1377.040 4.000 1377.640 ;
    END
  END bb_addr0[18]
  PIN bb_addr0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1406.960 4.000 1407.560 ;
    END
  END bb_addr0[19]
  PIN bb_addr0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 841.880 4.000 842.480 ;
    END
  END bb_addr0[1]
  PIN bb_addr0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1437.560 4.000 1438.160 ;
    END
  END bb_addr0[20]
  PIN bb_addr0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1468.160 4.000 1468.760 ;
    END
  END bb_addr0[21]
  PIN bb_addr0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1498.080 4.000 1498.680 ;
    END
  END bb_addr0[22]
  PIN bb_addr0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1528.680 4.000 1529.280 ;
    END
  END bb_addr0[23]
  PIN bb_addr0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1559.280 4.000 1559.880 ;
    END
  END bb_addr0[24]
  PIN bb_addr0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1589.880 4.000 1590.480 ;
    END
  END bb_addr0[25]
  PIN bb_addr0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1619.800 4.000 1620.400 ;
    END
  END bb_addr0[26]
  PIN bb_addr0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1650.400 4.000 1651.000 ;
    END
  END bb_addr0[27]
  PIN bb_addr0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1681.000 4.000 1681.600 ;
    END
  END bb_addr0[28]
  PIN bb_addr0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1710.920 4.000 1711.520 ;
    END
  END bb_addr0[29]
  PIN bb_addr0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 877.920 4.000 878.520 ;
    END
  END bb_addr0[2]
  PIN bb_addr0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1741.520 4.000 1742.120 ;
    END
  END bb_addr0[30]
  PIN bb_addr0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1772.120 4.000 1772.720 ;
    END
  END bb_addr0[31]
  PIN bb_addr0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 914.640 4.000 915.240 ;
    END
  END bb_addr0[3]
  PIN bb_addr0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 951.360 4.000 951.960 ;
    END
  END bb_addr0[4]
  PIN bb_addr0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 981.280 4.000 981.880 ;
    END
  END bb_addr0[5]
  PIN bb_addr0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1011.880 4.000 1012.480 ;
    END
  END bb_addr0[6]
  PIN bb_addr0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1042.480 4.000 1043.080 ;
    END
  END bb_addr0[7]
  PIN bb_addr0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1072.400 4.000 1073.000 ;
    END
  END bb_addr0[8]
  PIN bb_addr0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1103.000 4.000 1103.600 ;
    END
  END bb_addr0[9]
  PIN bb_addr1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 811.280 4.000 811.880 ;
    END
  END bb_addr1[0]
  PIN bb_addr1[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1139.720 4.000 1140.320 ;
    END
  END bb_addr1[10]
  PIN bb_addr1[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1169.640 4.000 1170.240 ;
    END
  END bb_addr1[11]
  PIN bb_addr1[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1200.240 4.000 1200.840 ;
    END
  END bb_addr1[12]
  PIN bb_addr1[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1230.840 4.000 1231.440 ;
    END
  END bb_addr1[13]
  PIN bb_addr1[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1261.440 4.000 1262.040 ;
    END
  END bb_addr1[14]
  PIN bb_addr1[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1291.360 4.000 1291.960 ;
    END
  END bb_addr1[15]
  PIN bb_addr1[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1321.960 4.000 1322.560 ;
    END
  END bb_addr1[16]
  PIN bb_addr1[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1352.560 4.000 1353.160 ;
    END
  END bb_addr1[17]
  PIN bb_addr1[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1382.480 4.000 1383.080 ;
    END
  END bb_addr1[18]
  PIN bb_addr1[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1413.080 4.000 1413.680 ;
    END
  END bb_addr1[19]
  PIN bb_addr1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 848.000 4.000 848.600 ;
    END
  END bb_addr1[1]
  PIN bb_addr1[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1443.680 4.000 1444.280 ;
    END
  END bb_addr1[20]
  PIN bb_addr1[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1474.280 4.000 1474.880 ;
    END
  END bb_addr1[21]
  PIN bb_addr1[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1504.200 4.000 1504.800 ;
    END
  END bb_addr1[22]
  PIN bb_addr1[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1534.800 4.000 1535.400 ;
    END
  END bb_addr1[23]
  PIN bb_addr1[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1565.400 4.000 1566.000 ;
    END
  END bb_addr1[24]
  PIN bb_addr1[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1595.320 4.000 1595.920 ;
    END
  END bb_addr1[25]
  PIN bb_addr1[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1625.920 4.000 1626.520 ;
    END
  END bb_addr1[26]
  PIN bb_addr1[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1656.520 4.000 1657.120 ;
    END
  END bb_addr1[27]
  PIN bb_addr1[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1687.120 4.000 1687.720 ;
    END
  END bb_addr1[28]
  PIN bb_addr1[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1717.040 4.000 1717.640 ;
    END
  END bb_addr1[29]
  PIN bb_addr1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 884.040 4.000 884.640 ;
    END
  END bb_addr1[2]
  PIN bb_addr1[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1747.640 4.000 1748.240 ;
    END
  END bb_addr1[30]
  PIN bb_addr1[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1778.240 4.000 1778.840 ;
    END
  END bb_addr1[31]
  PIN bb_addr1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 920.760 4.000 921.360 ;
    END
  END bb_addr1[3]
  PIN bb_addr1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 956.800 4.000 957.400 ;
    END
  END bb_addr1[4]
  PIN bb_addr1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 987.400 4.000 988.000 ;
    END
  END bb_addr1[5]
  PIN bb_addr1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1018.000 4.000 1018.600 ;
    END
  END bb_addr1[6]
  PIN bb_addr1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1048.600 4.000 1049.200 ;
    END
  END bb_addr1[7]
  PIN bb_addr1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1078.520 4.000 1079.120 ;
    END
  END bb_addr1[8]
  PIN bb_addr1[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1109.120 4.000 1109.720 ;
    END
  END bb_addr1[9]
  PIN bb_csb0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 786.800 4.000 787.400 ;
    END
  END bb_csb0
  PIN bb_csb1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 792.920 4.000 793.520 ;
    END
  END bb_csb1
  PIN bb_din0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 817.400 4.000 818.000 ;
    END
  END bb_din0[0]
  PIN bb_din0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1145.840 4.000 1146.440 ;
    END
  END bb_din0[10]
  PIN bb_din0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1175.760 4.000 1176.360 ;
    END
  END bb_din0[11]
  PIN bb_din0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1206.360 4.000 1206.960 ;
    END
  END bb_din0[12]
  PIN bb_din0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1236.960 4.000 1237.560 ;
    END
  END bb_din0[13]
  PIN bb_din0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1267.560 4.000 1268.160 ;
    END
  END bb_din0[14]
  PIN bb_din0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1297.480 4.000 1298.080 ;
    END
  END bb_din0[15]
  PIN bb_din0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1328.080 4.000 1328.680 ;
    END
  END bb_din0[16]
  PIN bb_din0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1358.680 4.000 1359.280 ;
    END
  END bb_din0[17]
  PIN bb_din0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1388.600 4.000 1389.200 ;
    END
  END bb_din0[18]
  PIN bb_din0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1419.200 4.000 1419.800 ;
    END
  END bb_din0[19]
  PIN bb_din0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 853.440 4.000 854.040 ;
    END
  END bb_din0[1]
  PIN bb_din0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1449.800 4.000 1450.400 ;
    END
  END bb_din0[20]
  PIN bb_din0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1480.400 4.000 1481.000 ;
    END
  END bb_din0[21]
  PIN bb_din0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1510.320 4.000 1510.920 ;
    END
  END bb_din0[22]
  PIN bb_din0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1540.920 4.000 1541.520 ;
    END
  END bb_din0[23]
  PIN bb_din0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1571.520 4.000 1572.120 ;
    END
  END bb_din0[24]
  PIN bb_din0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1601.440 4.000 1602.040 ;
    END
  END bb_din0[25]
  PIN bb_din0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1632.040 4.000 1632.640 ;
    END
  END bb_din0[26]
  PIN bb_din0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1662.640 4.000 1663.240 ;
    END
  END bb_din0[27]
  PIN bb_din0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1693.240 4.000 1693.840 ;
    END
  END bb_din0[28]
  PIN bb_din0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1723.160 4.000 1723.760 ;
    END
  END bb_din0[29]
  PIN bb_din0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 890.160 4.000 890.760 ;
    END
  END bb_din0[2]
  PIN bb_din0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1753.760 4.000 1754.360 ;
    END
  END bb_din0[30]
  PIN bb_din0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1784.360 4.000 1784.960 ;
    END
  END bb_din0[31]
  PIN bb_din0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 926.880 4.000 927.480 ;
    END
  END bb_din0[3]
  PIN bb_din0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 962.920 4.000 963.520 ;
    END
  END bb_din0[4]
  PIN bb_din0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 993.520 4.000 994.120 ;
    END
  END bb_din0[5]
  PIN bb_din0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1024.120 4.000 1024.720 ;
    END
  END bb_din0[6]
  PIN bb_din0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1054.720 4.000 1055.320 ;
    END
  END bb_din0[7]
  PIN bb_din0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1084.640 4.000 1085.240 ;
    END
  END bb_din0[8]
  PIN bb_din0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1115.240 4.000 1115.840 ;
    END
  END bb_din0[9]
  PIN bb_dout0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 823.520 4.000 824.120 ;
    END
  END bb_dout0[0]
  PIN bb_dout0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1151.960 4.000 1152.560 ;
    END
  END bb_dout0[10]
  PIN bb_dout0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1181.880 4.000 1182.480 ;
    END
  END bb_dout0[11]
  PIN bb_dout0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1212.480 4.000 1213.080 ;
    END
  END bb_dout0[12]
  PIN bb_dout0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1243.080 4.000 1243.680 ;
    END
  END bb_dout0[13]
  PIN bb_dout0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1273.000 4.000 1273.600 ;
    END
  END bb_dout0[14]
  PIN bb_dout0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1303.600 4.000 1304.200 ;
    END
  END bb_dout0[15]
  PIN bb_dout0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1334.200 4.000 1334.800 ;
    END
  END bb_dout0[16]
  PIN bb_dout0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1364.800 4.000 1365.400 ;
    END
  END bb_dout0[17]
  PIN bb_dout0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1394.720 4.000 1395.320 ;
    END
  END bb_dout0[18]
  PIN bb_dout0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1425.320 4.000 1425.920 ;
    END
  END bb_dout0[19]
  PIN bb_dout0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 859.560 4.000 860.160 ;
    END
  END bb_dout0[1]
  PIN bb_dout0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1455.920 4.000 1456.520 ;
    END
  END bb_dout0[20]
  PIN bb_dout0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1485.840 4.000 1486.440 ;
    END
  END bb_dout0[21]
  PIN bb_dout0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1516.440 4.000 1517.040 ;
    END
  END bb_dout0[22]
  PIN bb_dout0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1547.040 4.000 1547.640 ;
    END
  END bb_dout0[23]
  PIN bb_dout0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1577.640 4.000 1578.240 ;
    END
  END bb_dout0[24]
  PIN bb_dout0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1607.560 4.000 1608.160 ;
    END
  END bb_dout0[25]
  PIN bb_dout0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1638.160 4.000 1638.760 ;
    END
  END bb_dout0[26]
  PIN bb_dout0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1668.760 4.000 1669.360 ;
    END
  END bb_dout0[27]
  PIN bb_dout0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1698.680 4.000 1699.280 ;
    END
  END bb_dout0[28]
  PIN bb_dout0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1729.280 4.000 1729.880 ;
    END
  END bb_dout0[29]
  PIN bb_dout0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 896.280 4.000 896.880 ;
    END
  END bb_dout0[2]
  PIN bb_dout0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1759.880 4.000 1760.480 ;
    END
  END bb_dout0[30]
  PIN bb_dout0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1790.480 4.000 1791.080 ;
    END
  END bb_dout0[31]
  PIN bb_dout0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 933.000 4.000 933.600 ;
    END
  END bb_dout0[3]
  PIN bb_dout0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 969.040 4.000 969.640 ;
    END
  END bb_dout0[4]
  PIN bb_dout0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 999.640 4.000 1000.240 ;
    END
  END bb_dout0[5]
  PIN bb_dout0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1030.240 4.000 1030.840 ;
    END
  END bb_dout0[6]
  PIN bb_dout0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1060.840 4.000 1061.440 ;
    END
  END bb_dout0[7]
  PIN bb_dout0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1090.760 4.000 1091.360 ;
    END
  END bb_dout0[8]
  PIN bb_dout0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1121.360 4.000 1121.960 ;
    END
  END bb_dout0[9]
  PIN bb_dout1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 829.640 4.000 830.240 ;
    END
  END bb_dout1[0]
  PIN bb_dout1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1158.080 4.000 1158.680 ;
    END
  END bb_dout1[10]
  PIN bb_dout1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1188.000 4.000 1188.600 ;
    END
  END bb_dout1[11]
  PIN bb_dout1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1218.600 4.000 1219.200 ;
    END
  END bb_dout1[12]
  PIN bb_dout1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1249.200 4.000 1249.800 ;
    END
  END bb_dout1[13]
  PIN bb_dout1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1279.120 4.000 1279.720 ;
    END
  END bb_dout1[14]
  PIN bb_dout1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1309.720 4.000 1310.320 ;
    END
  END bb_dout1[15]
  PIN bb_dout1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1340.320 4.000 1340.920 ;
    END
  END bb_dout1[16]
  PIN bb_dout1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1370.920 4.000 1371.520 ;
    END
  END bb_dout1[17]
  PIN bb_dout1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1400.840 4.000 1401.440 ;
    END
  END bb_dout1[18]
  PIN bb_dout1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1431.440 4.000 1432.040 ;
    END
  END bb_dout1[19]
  PIN bb_dout1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 865.680 4.000 866.280 ;
    END
  END bb_dout1[1]
  PIN bb_dout1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1462.040 4.000 1462.640 ;
    END
  END bb_dout1[20]
  PIN bb_dout1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1491.960 4.000 1492.560 ;
    END
  END bb_dout1[21]
  PIN bb_dout1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1522.560 4.000 1523.160 ;
    END
  END bb_dout1[22]
  PIN bb_dout1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1553.160 4.000 1553.760 ;
    END
  END bb_dout1[23]
  PIN bb_dout1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1583.760 4.000 1584.360 ;
    END
  END bb_dout1[24]
  PIN bb_dout1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1613.680 4.000 1614.280 ;
    END
  END bb_dout1[25]
  PIN bb_dout1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1644.280 4.000 1644.880 ;
    END
  END bb_dout1[26]
  PIN bb_dout1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1674.880 4.000 1675.480 ;
    END
  END bb_dout1[27]
  PIN bb_dout1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1704.800 4.000 1705.400 ;
    END
  END bb_dout1[28]
  PIN bb_dout1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1735.400 4.000 1736.000 ;
    END
  END bb_dout1[29]
  PIN bb_dout1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 902.400 4.000 903.000 ;
    END
  END bb_dout1[2]
  PIN bb_dout1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1766.000 4.000 1766.600 ;
    END
  END bb_dout1[30]
  PIN bb_dout1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1796.600 4.000 1797.200 ;
    END
  END bb_dout1[31]
  PIN bb_dout1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 939.120 4.000 939.720 ;
    END
  END bb_dout1[3]
  PIN bb_dout1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 975.160 4.000 975.760 ;
    END
  END bb_dout1[4]
  PIN bb_dout1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1005.760 4.000 1006.360 ;
    END
  END bb_dout1[5]
  PIN bb_dout1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1036.360 4.000 1036.960 ;
    END
  END bb_dout1[6]
  PIN bb_dout1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1066.280 4.000 1066.880 ;
    END
  END bb_dout1[7]
  PIN bb_dout1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1096.880 4.000 1097.480 ;
    END
  END bb_dout1[8]
  PIN bb_dout1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1127.480 4.000 1128.080 ;
    END
  END bb_dout1[9]
  PIN bb_web0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 799.040 4.000 799.640 ;
    END
  END bb_web0
  PIN bb_wmask0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 835.760 4.000 836.360 ;
    END
  END bb_wmask0[0]
  PIN bb_wmask0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 871.800 4.000 872.400 ;
    END
  END bb_wmask0[1]
  PIN bb_wmask0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 908.520 4.000 909.120 ;
    END
  END bb_wmask0[2]
  PIN bb_wmask0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 945.240 4.000 945.840 ;
    END
  END bb_wmask0[3]
  PIN clk_g
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.910 0.000 8.190 4.000 ;
    END
  END clk_g
  PIN io_gecerli
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.850 0.000 72.130 4.000 ;
    END
  END io_gecerli
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.490 0.000 87.770 4.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 407.650 0.000 407.930 4.000 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 439.850 0.000 440.130 4.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 471.590 0.000 471.870 4.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 503.790 0.000 504.070 4.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 535.530 0.000 535.810 4.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 567.730 0.000 568.010 4.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.930 0.000 600.210 4.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 631.670 0.000 631.950 4.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 663.870 0.000 664.150 4.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 695.610 0.000 695.890 4.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.690 0.000 119.970 4.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 727.810 0.000 728.090 4.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 759.550 0.000 759.830 4.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 791.750 0.000 792.030 4.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 823.950 0.000 824.230 4.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 855.690 0.000 855.970 4.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 887.890 0.000 888.170 4.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 919.630 0.000 919.910 4.000 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 951.830 0.000 952.110 4.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 983.570 0.000 983.850 4.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1015.770 0.000 1016.050 4.000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.890 0.000 152.170 4.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1047.970 0.000 1048.250 4.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1079.710 0.000 1079.990 4.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1111.910 0.000 1112.190 4.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1128.010 0.000 1128.290 4.000 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1143.650 0.000 1143.930 4.000 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1159.750 0.000 1160.030 4.000 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1175.850 0.000 1176.130 4.000 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1191.950 0.000 1192.230 4.000 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.630 0.000 183.910 4.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.830 0.000 216.110 4.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.570 0.000 247.850 4.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.770 0.000 280.050 4.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.510 0.000 311.790 4.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 343.710 0.000 343.990 4.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 375.910 0.000 376.190 4.000 ;
    END
  END io_oeb[9]
  PIN io_ps[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.590 0.000 103.870 4.000 ;
    END
  END io_ps[0]
  PIN io_ps[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 423.750 0.000 424.030 4.000 ;
    END
  END io_ps[10]
  PIN io_ps[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 455.950 0.000 456.230 4.000 ;
    END
  END io_ps[11]
  PIN io_ps[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 487.690 0.000 487.970 4.000 ;
    END
  END io_ps[12]
  PIN io_ps[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 519.890 0.000 520.170 4.000 ;
    END
  END io_ps[13]
  PIN io_ps[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 551.630 0.000 551.910 4.000 ;
    END
  END io_ps[14]
  PIN io_ps[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 583.830 0.000 584.110 4.000 ;
    END
  END io_ps[15]
  PIN io_ps[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 615.570 0.000 615.850 4.000 ;
    END
  END io_ps[16]
  PIN io_ps[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 647.770 0.000 648.050 4.000 ;
    END
  END io_ps[17]
  PIN io_ps[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 679.970 0.000 680.250 4.000 ;
    END
  END io_ps[18]
  PIN io_ps[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 711.710 0.000 711.990 4.000 ;
    END
  END io_ps[19]
  PIN io_ps[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.790 0.000 136.070 4.000 ;
    END
  END io_ps[1]
  PIN io_ps[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 743.910 0.000 744.190 4.000 ;
    END
  END io_ps[20]
  PIN io_ps[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 775.650 0.000 775.930 4.000 ;
    END
  END io_ps[21]
  PIN io_ps[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 807.850 0.000 808.130 4.000 ;
    END
  END io_ps[22]
  PIN io_ps[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 839.590 0.000 839.870 4.000 ;
    END
  END io_ps[23]
  PIN io_ps[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 871.790 0.000 872.070 4.000 ;
    END
  END io_ps[24]
  PIN io_ps[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 903.990 0.000 904.270 4.000 ;
    END
  END io_ps[25]
  PIN io_ps[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 935.730 0.000 936.010 4.000 ;
    END
  END io_ps[26]
  PIN io_ps[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 967.930 0.000 968.210 4.000 ;
    END
  END io_ps[27]
  PIN io_ps[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 999.670 0.000 999.950 4.000 ;
    END
  END io_ps[28]
  PIN io_ps[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1031.870 0.000 1032.150 4.000 ;
    END
  END io_ps[29]
  PIN io_ps[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 0.000 167.810 4.000 ;
    END
  END io_ps[2]
  PIN io_ps[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1063.610 0.000 1063.890 4.000 ;
    END
  END io_ps[30]
  PIN io_ps[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1095.810 0.000 1096.090 4.000 ;
    END
  END io_ps[31]
  PIN io_ps[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.730 0.000 200.010 4.000 ;
    END
  END io_ps[3]
  PIN io_ps[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.930 0.000 232.210 4.000 ;
    END
  END io_ps[4]
  PIN io_ps[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.670 0.000 263.950 4.000 ;
    END
  END io_ps[5]
  PIN io_ps[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 295.870 0.000 296.150 4.000 ;
    END
  END io_ps[6]
  PIN io_ps[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 327.610 0.000 327.890 4.000 ;
    END
  END io_ps[7]
  PIN io_ps[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 359.810 0.000 360.090 4.000 ;
    END
  END io_ps[8]
  PIN io_ps[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 391.550 0.000 391.830 4.000 ;
    END
  END io_ps[9]
  PIN rst_g
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.550 0.000 23.830 4.000 ;
    END
  END rst_g
  PIN rx
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.750 0.000 56.030 4.000 ;
    END
  END rx
  PIN tx
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.650 0.000 39.930 4.000 ;
    END
  END tx
  PIN vb_addr0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END vb_addr0[0]
  PIN vb_addr0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 348.880 4.000 349.480 ;
    END
  END vb_addr0[10]
  PIN vb_addr0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 379.480 4.000 380.080 ;
    END
  END vb_addr0[11]
  PIN vb_addr0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 410.080 4.000 410.680 ;
    END
  END vb_addr0[12]
  PIN vb_addr0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.160 4.000 57.760 ;
    END
  END vb_addr0[1]
  PIN vb_addr0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.880 4.000 94.480 ;
    END
  END vb_addr0[2]
  PIN vb_addr0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.920 4.000 130.520 ;
    END
  END vb_addr0[3]
  PIN vb_addr0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 166.640 4.000 167.240 ;
    END
  END vb_addr0[4]
  PIN vb_addr0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 197.240 4.000 197.840 ;
    END
  END vb_addr0[5]
  PIN vb_addr0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.160 4.000 227.760 ;
    END
  END vb_addr0[6]
  PIN vb_addr0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 257.760 4.000 258.360 ;
    END
  END vb_addr0[7]
  PIN vb_addr0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 288.360 4.000 288.960 ;
    END
  END vb_addr0[8]
  PIN vb_addr0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 318.960 4.000 319.560 ;
    END
  END vb_addr0[9]
  PIN vb_addr1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 26.560 4.000 27.160 ;
    END
  END vb_addr1[0]
  PIN vb_addr1[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 355.000 4.000 355.600 ;
    END
  END vb_addr1[10]
  PIN vb_addr1[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 385.600 4.000 386.200 ;
    END
  END vb_addr1[11]
  PIN vb_addr1[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 416.200 4.000 416.800 ;
    END
  END vb_addr1[12]
  PIN vb_addr1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.280 4.000 63.880 ;
    END
  END vb_addr1[1]
  PIN vb_addr1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.000 4.000 100.600 ;
    END
  END vb_addr1[2]
  PIN vb_addr1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.040 4.000 136.640 ;
    END
  END vb_addr1[3]
  PIN vb_addr1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 172.760 4.000 173.360 ;
    END
  END vb_addr1[4]
  PIN vb_addr1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 203.360 4.000 203.960 ;
    END
  END vb_addr1[5]
  PIN vb_addr1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 233.280 4.000 233.880 ;
    END
  END vb_addr1[6]
  PIN vb_addr1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 263.880 4.000 264.480 ;
    END
  END vb_addr1[7]
  PIN vb_addr1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 294.480 4.000 295.080 ;
    END
  END vb_addr1[8]
  PIN vb_addr1[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 324.400 4.000 325.000 ;
    END
  END vb_addr1[9]
  PIN vb_csb0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.760 4.000 3.360 ;
    END
  END vb_csb0
  PIN vb_csb1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.200 4.000 8.800 ;
    END
  END vb_csb1
  PIN vb_din0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.680 4.000 33.280 ;
    END
  END vb_din0[0]
  PIN vb_din0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 361.120 4.000 361.720 ;
    END
  END vb_din0[10]
  PIN vb_din0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 391.720 4.000 392.320 ;
    END
  END vb_din0[11]
  PIN vb_din0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 422.320 4.000 422.920 ;
    END
  END vb_din0[12]
  PIN vb_din0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 440.000 4.000 440.600 ;
    END
  END vb_din0[13]
  PIN vb_din0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 458.360 4.000 458.960 ;
    END
  END vb_din0[14]
  PIN vb_din0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 476.720 4.000 477.320 ;
    END
  END vb_din0[15]
  PIN vb_din0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 495.080 4.000 495.680 ;
    END
  END vb_din0[16]
  PIN vb_din0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 513.440 4.000 514.040 ;
    END
  END vb_din0[17]
  PIN vb_din0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 531.800 4.000 532.400 ;
    END
  END vb_din0[18]
  PIN vb_din0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 549.480 4.000 550.080 ;
    END
  END vb_din0[19]
  PIN vb_din0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 69.400 4.000 70.000 ;
    END
  END vb_din0[1]
  PIN vb_din0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 567.840 4.000 568.440 ;
    END
  END vb_din0[20]
  PIN vb_din0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 586.200 4.000 586.800 ;
    END
  END vb_din0[21]
  PIN vb_din0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 604.560 4.000 605.160 ;
    END
  END vb_din0[22]
  PIN vb_din0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 622.920 4.000 623.520 ;
    END
  END vb_din0[23]
  PIN vb_din0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 640.600 4.000 641.200 ;
    END
  END vb_din0[24]
  PIN vb_din0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 658.960 4.000 659.560 ;
    END
  END vb_din0[25]
  PIN vb_din0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 677.320 4.000 677.920 ;
    END
  END vb_din0[26]
  PIN vb_din0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 695.680 4.000 696.280 ;
    END
  END vb_din0[27]
  PIN vb_din0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 714.040 4.000 714.640 ;
    END
  END vb_din0[28]
  PIN vb_din0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 732.400 4.000 733.000 ;
    END
  END vb_din0[29]
  PIN vb_din0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.120 4.000 106.720 ;
    END
  END vb_din0[2]
  PIN vb_din0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 750.080 4.000 750.680 ;
    END
  END vb_din0[30]
  PIN vb_din0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 768.440 4.000 769.040 ;
    END
  END vb_din0[31]
  PIN vb_din0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.160 4.000 142.760 ;
    END
  END vb_din0[3]
  PIN vb_din0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 178.880 4.000 179.480 ;
    END
  END vb_din0[4]
  PIN vb_din0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 209.480 4.000 210.080 ;
    END
  END vb_din0[5]
  PIN vb_din0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 239.400 4.000 240.000 ;
    END
  END vb_din0[6]
  PIN vb_din0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 270.000 4.000 270.600 ;
    END
  END vb_din0[7]
  PIN vb_din0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 300.600 4.000 301.200 ;
    END
  END vb_din0[8]
  PIN vb_din0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 330.520 4.000 331.120 ;
    END
  END vb_din0[9]
  PIN vb_dout0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.800 4.000 39.400 ;
    END
  END vb_dout0[0]
  PIN vb_dout0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 367.240 4.000 367.840 ;
    END
  END vb_dout0[10]
  PIN vb_dout0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 397.840 4.000 398.440 ;
    END
  END vb_dout0[11]
  PIN vb_dout0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 427.760 4.000 428.360 ;
    END
  END vb_dout0[12]
  PIN vb_dout0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 446.120 4.000 446.720 ;
    END
  END vb_dout0[13]
  PIN vb_dout0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 464.480 4.000 465.080 ;
    END
  END vb_dout0[14]
  PIN vb_dout0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 482.840 4.000 483.440 ;
    END
  END vb_dout0[15]
  PIN vb_dout0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 501.200 4.000 501.800 ;
    END
  END vb_dout0[16]
  PIN vb_dout0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 519.560 4.000 520.160 ;
    END
  END vb_dout0[17]
  PIN vb_dout0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 537.240 4.000 537.840 ;
    END
  END vb_dout0[18]
  PIN vb_dout0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 555.600 4.000 556.200 ;
    END
  END vb_dout0[19]
  PIN vb_dout0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 75.520 4.000 76.120 ;
    END
  END vb_dout0[1]
  PIN vb_dout0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 573.960 4.000 574.560 ;
    END
  END vb_dout0[20]
  PIN vb_dout0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 592.320 4.000 592.920 ;
    END
  END vb_dout0[21]
  PIN vb_dout0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 610.680 4.000 611.280 ;
    END
  END vb_dout0[22]
  PIN vb_dout0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 629.040 4.000 629.640 ;
    END
  END vb_dout0[23]
  PIN vb_dout0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 646.720 4.000 647.320 ;
    END
  END vb_dout0[24]
  PIN vb_dout0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 665.080 4.000 665.680 ;
    END
  END vb_dout0[25]
  PIN vb_dout0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 683.440 4.000 684.040 ;
    END
  END vb_dout0[26]
  PIN vb_dout0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 701.800 4.000 702.400 ;
    END
  END vb_dout0[27]
  PIN vb_dout0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 720.160 4.000 720.760 ;
    END
  END vb_dout0[28]
  PIN vb_dout0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 738.520 4.000 739.120 ;
    END
  END vb_dout0[29]
  PIN vb_dout0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 111.560 4.000 112.160 ;
    END
  END vb_dout0[2]
  PIN vb_dout0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 756.200 4.000 756.800 ;
    END
  END vb_dout0[30]
  PIN vb_dout0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 774.560 4.000 775.160 ;
    END
  END vb_dout0[31]
  PIN vb_dout0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 148.280 4.000 148.880 ;
    END
  END vb_dout0[3]
  PIN vb_dout0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 185.000 4.000 185.600 ;
    END
  END vb_dout0[4]
  PIN vb_dout0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.920 4.000 215.520 ;
    END
  END vb_dout0[5]
  PIN vb_dout0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 245.520 4.000 246.120 ;
    END
  END vb_dout0[6]
  PIN vb_dout0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 276.120 4.000 276.720 ;
    END
  END vb_dout0[7]
  PIN vb_dout0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 306.720 4.000 307.320 ;
    END
  END vb_dout0[8]
  PIN vb_dout0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 336.640 4.000 337.240 ;
    END
  END vb_dout0[9]
  PIN vb_dout1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.920 4.000 45.520 ;
    END
  END vb_dout1[0]
  PIN vb_dout1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 373.360 4.000 373.960 ;
    END
  END vb_dout1[10]
  PIN vb_dout1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 403.960 4.000 404.560 ;
    END
  END vb_dout1[11]
  PIN vb_dout1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 433.880 4.000 434.480 ;
    END
  END vb_dout1[12]
  PIN vb_dout1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 452.240 4.000 452.840 ;
    END
  END vb_dout1[13]
  PIN vb_dout1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 470.600 4.000 471.200 ;
    END
  END vb_dout1[14]
  PIN vb_dout1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 488.960 4.000 489.560 ;
    END
  END vb_dout1[15]
  PIN vb_dout1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 507.320 4.000 507.920 ;
    END
  END vb_dout1[16]
  PIN vb_dout1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 525.680 4.000 526.280 ;
    END
  END vb_dout1[17]
  PIN vb_dout1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 543.360 4.000 543.960 ;
    END
  END vb_dout1[18]
  PIN vb_dout1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 561.720 4.000 562.320 ;
    END
  END vb_dout1[19]
  PIN vb_dout1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END vb_dout1[1]
  PIN vb_dout1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 580.080 4.000 580.680 ;
    END
  END vb_dout1[20]
  PIN vb_dout1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 598.440 4.000 599.040 ;
    END
  END vb_dout1[21]
  PIN vb_dout1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 616.800 4.000 617.400 ;
    END
  END vb_dout1[22]
  PIN vb_dout1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 635.160 4.000 635.760 ;
    END
  END vb_dout1[23]
  PIN vb_dout1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 652.840 4.000 653.440 ;
    END
  END vb_dout1[24]
  PIN vb_dout1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 671.200 4.000 671.800 ;
    END
  END vb_dout1[25]
  PIN vb_dout1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 689.560 4.000 690.160 ;
    END
  END vb_dout1[26]
  PIN vb_dout1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 707.920 4.000 708.520 ;
    END
  END vb_dout1[27]
  PIN vb_dout1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 726.280 4.000 726.880 ;
    END
  END vb_dout1[28]
  PIN vb_dout1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 743.960 4.000 744.560 ;
    END
  END vb_dout1[29]
  PIN vb_dout1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.680 4.000 118.280 ;
    END
  END vb_dout1[2]
  PIN vb_dout1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 762.320 4.000 762.920 ;
    END
  END vb_dout1[30]
  PIN vb_dout1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 780.680 4.000 781.280 ;
    END
  END vb_dout1[31]
  PIN vb_dout1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 154.400 4.000 155.000 ;
    END
  END vb_dout1[3]
  PIN vb_dout1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 191.120 4.000 191.720 ;
    END
  END vb_dout1[4]
  PIN vb_dout1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 221.040 4.000 221.640 ;
    END
  END vb_dout1[5]
  PIN vb_dout1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 251.640 4.000 252.240 ;
    END
  END vb_dout1[6]
  PIN vb_dout1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 282.240 4.000 282.840 ;
    END
  END vb_dout1[7]
  PIN vb_dout1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 312.840 4.000 313.440 ;
    END
  END vb_dout1[8]
  PIN vb_dout1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 342.760 4.000 343.360 ;
    END
  END vb_dout1[9]
  PIN vb_web0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 14.320 4.000 14.920 ;
    END
  END vb_web0
  PIN vb_wmask0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 4.000 51.640 ;
    END
  END vb_wmask0[0]
  PIN vb_wmask0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 87.760 4.000 88.360 ;
    END
  END vb_wmask0[1]
  PIN vb_wmask0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 123.800 4.000 124.400 ;
    END
  END vb_wmask0[2]
  PIN vb_wmask0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 160.520 4.000 161.120 ;
    END
  END vb_wmask0[3]
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1787.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 1787.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 1787.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 1787.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 1787.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 1787.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 1787.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 1787.280 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 1787.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 1787.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 1787.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 1787.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 1787.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 1787.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 1787.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 1787.280 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 1194.160 1787.125 ;
      LAYER met1 ;
        RECT 3.750 10.640 1194.160 1787.280 ;
      LAYER met2 ;
        RECT 3.780 4.280 1192.220 1797.085 ;
        RECT 3.780 2.875 7.630 4.280 ;
        RECT 8.470 2.875 23.270 4.280 ;
        RECT 24.110 2.875 39.370 4.280 ;
        RECT 40.210 2.875 55.470 4.280 ;
        RECT 56.310 2.875 71.570 4.280 ;
        RECT 72.410 2.875 87.210 4.280 ;
        RECT 88.050 2.875 103.310 4.280 ;
        RECT 104.150 2.875 119.410 4.280 ;
        RECT 120.250 2.875 135.510 4.280 ;
        RECT 136.350 2.875 151.610 4.280 ;
        RECT 152.450 2.875 167.250 4.280 ;
        RECT 168.090 2.875 183.350 4.280 ;
        RECT 184.190 2.875 199.450 4.280 ;
        RECT 200.290 2.875 215.550 4.280 ;
        RECT 216.390 2.875 231.650 4.280 ;
        RECT 232.490 2.875 247.290 4.280 ;
        RECT 248.130 2.875 263.390 4.280 ;
        RECT 264.230 2.875 279.490 4.280 ;
        RECT 280.330 2.875 295.590 4.280 ;
        RECT 296.430 2.875 311.230 4.280 ;
        RECT 312.070 2.875 327.330 4.280 ;
        RECT 328.170 2.875 343.430 4.280 ;
        RECT 344.270 2.875 359.530 4.280 ;
        RECT 360.370 2.875 375.630 4.280 ;
        RECT 376.470 2.875 391.270 4.280 ;
        RECT 392.110 2.875 407.370 4.280 ;
        RECT 408.210 2.875 423.470 4.280 ;
        RECT 424.310 2.875 439.570 4.280 ;
        RECT 440.410 2.875 455.670 4.280 ;
        RECT 456.510 2.875 471.310 4.280 ;
        RECT 472.150 2.875 487.410 4.280 ;
        RECT 488.250 2.875 503.510 4.280 ;
        RECT 504.350 2.875 519.610 4.280 ;
        RECT 520.450 2.875 535.250 4.280 ;
        RECT 536.090 2.875 551.350 4.280 ;
        RECT 552.190 2.875 567.450 4.280 ;
        RECT 568.290 2.875 583.550 4.280 ;
        RECT 584.390 2.875 599.650 4.280 ;
        RECT 600.490 2.875 615.290 4.280 ;
        RECT 616.130 2.875 631.390 4.280 ;
        RECT 632.230 2.875 647.490 4.280 ;
        RECT 648.330 2.875 663.590 4.280 ;
        RECT 664.430 2.875 679.690 4.280 ;
        RECT 680.530 2.875 695.330 4.280 ;
        RECT 696.170 2.875 711.430 4.280 ;
        RECT 712.270 2.875 727.530 4.280 ;
        RECT 728.370 2.875 743.630 4.280 ;
        RECT 744.470 2.875 759.270 4.280 ;
        RECT 760.110 2.875 775.370 4.280 ;
        RECT 776.210 2.875 791.470 4.280 ;
        RECT 792.310 2.875 807.570 4.280 ;
        RECT 808.410 2.875 823.670 4.280 ;
        RECT 824.510 2.875 839.310 4.280 ;
        RECT 840.150 2.875 855.410 4.280 ;
        RECT 856.250 2.875 871.510 4.280 ;
        RECT 872.350 2.875 887.610 4.280 ;
        RECT 888.450 2.875 903.710 4.280 ;
        RECT 904.550 2.875 919.350 4.280 ;
        RECT 920.190 2.875 935.450 4.280 ;
        RECT 936.290 2.875 951.550 4.280 ;
        RECT 952.390 2.875 967.650 4.280 ;
        RECT 968.490 2.875 983.290 4.280 ;
        RECT 984.130 2.875 999.390 4.280 ;
        RECT 1000.230 2.875 1015.490 4.280 ;
        RECT 1016.330 2.875 1031.590 4.280 ;
        RECT 1032.430 2.875 1047.690 4.280 ;
        RECT 1048.530 2.875 1063.330 4.280 ;
        RECT 1064.170 2.875 1079.430 4.280 ;
        RECT 1080.270 2.875 1095.530 4.280 ;
        RECT 1096.370 2.875 1111.630 4.280 ;
        RECT 1112.470 2.875 1127.730 4.280 ;
        RECT 1128.570 2.875 1143.370 4.280 ;
        RECT 1144.210 2.875 1159.470 4.280 ;
        RECT 1160.310 2.875 1175.570 4.280 ;
        RECT 1176.410 2.875 1191.670 4.280 ;
      LAYER met3 ;
        RECT 4.400 1796.200 1174.640 1797.065 ;
        RECT 4.000 1791.480 1174.640 1796.200 ;
        RECT 4.400 1790.080 1174.640 1791.480 ;
        RECT 4.000 1785.360 1174.640 1790.080 ;
        RECT 4.400 1783.960 1174.640 1785.360 ;
        RECT 4.000 1779.240 1174.640 1783.960 ;
        RECT 4.400 1777.840 1174.640 1779.240 ;
        RECT 4.000 1773.120 1174.640 1777.840 ;
        RECT 4.400 1771.720 1174.640 1773.120 ;
        RECT 4.000 1767.000 1174.640 1771.720 ;
        RECT 4.400 1765.600 1174.640 1767.000 ;
        RECT 4.000 1760.880 1174.640 1765.600 ;
        RECT 4.400 1759.480 1174.640 1760.880 ;
        RECT 4.000 1754.760 1174.640 1759.480 ;
        RECT 4.400 1753.360 1174.640 1754.760 ;
        RECT 4.000 1748.640 1174.640 1753.360 ;
        RECT 4.400 1747.240 1174.640 1748.640 ;
        RECT 4.000 1742.520 1174.640 1747.240 ;
        RECT 4.400 1741.120 1174.640 1742.520 ;
        RECT 4.000 1736.400 1174.640 1741.120 ;
        RECT 4.400 1735.000 1174.640 1736.400 ;
        RECT 4.000 1730.280 1174.640 1735.000 ;
        RECT 4.400 1728.880 1174.640 1730.280 ;
        RECT 4.000 1724.160 1174.640 1728.880 ;
        RECT 4.400 1722.760 1174.640 1724.160 ;
        RECT 4.000 1718.040 1174.640 1722.760 ;
        RECT 4.400 1716.640 1174.640 1718.040 ;
        RECT 4.000 1711.920 1174.640 1716.640 ;
        RECT 4.400 1710.520 1174.640 1711.920 ;
        RECT 4.000 1705.800 1174.640 1710.520 ;
        RECT 4.400 1704.400 1174.640 1705.800 ;
        RECT 4.000 1699.680 1174.640 1704.400 ;
        RECT 4.400 1698.280 1174.640 1699.680 ;
        RECT 4.000 1694.240 1174.640 1698.280 ;
        RECT 4.400 1692.840 1174.640 1694.240 ;
        RECT 4.000 1688.120 1174.640 1692.840 ;
        RECT 4.400 1686.720 1174.640 1688.120 ;
        RECT 4.000 1682.000 1174.640 1686.720 ;
        RECT 4.400 1680.600 1174.640 1682.000 ;
        RECT 4.000 1675.880 1174.640 1680.600 ;
        RECT 4.400 1674.480 1174.640 1675.880 ;
        RECT 4.000 1669.760 1174.640 1674.480 ;
        RECT 4.400 1668.360 1174.640 1669.760 ;
        RECT 4.000 1663.640 1174.640 1668.360 ;
        RECT 4.400 1662.240 1174.640 1663.640 ;
        RECT 4.000 1657.520 1174.640 1662.240 ;
        RECT 4.400 1656.120 1174.640 1657.520 ;
        RECT 4.000 1651.400 1174.640 1656.120 ;
        RECT 4.400 1650.000 1174.640 1651.400 ;
        RECT 4.000 1645.280 1174.640 1650.000 ;
        RECT 4.400 1643.880 1174.640 1645.280 ;
        RECT 4.000 1639.160 1174.640 1643.880 ;
        RECT 4.400 1637.760 1174.640 1639.160 ;
        RECT 4.000 1633.040 1174.640 1637.760 ;
        RECT 4.400 1631.640 1174.640 1633.040 ;
        RECT 4.000 1626.920 1174.640 1631.640 ;
        RECT 4.400 1625.520 1174.640 1626.920 ;
        RECT 4.000 1620.800 1174.640 1625.520 ;
        RECT 4.400 1619.400 1174.640 1620.800 ;
        RECT 4.000 1614.680 1174.640 1619.400 ;
        RECT 4.400 1613.280 1174.640 1614.680 ;
        RECT 4.000 1608.560 1174.640 1613.280 ;
        RECT 4.400 1607.160 1174.640 1608.560 ;
        RECT 4.000 1602.440 1174.640 1607.160 ;
        RECT 4.400 1601.040 1174.640 1602.440 ;
        RECT 4.000 1596.320 1174.640 1601.040 ;
        RECT 4.400 1594.920 1174.640 1596.320 ;
        RECT 4.000 1590.880 1174.640 1594.920 ;
        RECT 4.400 1589.480 1174.640 1590.880 ;
        RECT 4.000 1584.760 1174.640 1589.480 ;
        RECT 4.400 1583.360 1174.640 1584.760 ;
        RECT 4.000 1578.640 1174.640 1583.360 ;
        RECT 4.400 1577.240 1174.640 1578.640 ;
        RECT 4.000 1572.520 1174.640 1577.240 ;
        RECT 4.400 1571.120 1174.640 1572.520 ;
        RECT 4.000 1566.400 1174.640 1571.120 ;
        RECT 4.400 1565.000 1174.640 1566.400 ;
        RECT 4.000 1560.280 1174.640 1565.000 ;
        RECT 4.400 1558.880 1174.640 1560.280 ;
        RECT 4.000 1554.160 1174.640 1558.880 ;
        RECT 4.400 1552.760 1174.640 1554.160 ;
        RECT 4.000 1548.040 1174.640 1552.760 ;
        RECT 4.400 1546.640 1174.640 1548.040 ;
        RECT 4.000 1541.920 1174.640 1546.640 ;
        RECT 4.400 1540.520 1174.640 1541.920 ;
        RECT 4.000 1535.800 1174.640 1540.520 ;
        RECT 4.400 1534.400 1174.640 1535.800 ;
        RECT 4.000 1529.680 1174.640 1534.400 ;
        RECT 4.400 1528.280 1174.640 1529.680 ;
        RECT 4.000 1523.560 1174.640 1528.280 ;
        RECT 4.400 1522.160 1174.640 1523.560 ;
        RECT 4.000 1517.440 1174.640 1522.160 ;
        RECT 4.400 1516.040 1174.640 1517.440 ;
        RECT 4.000 1511.320 1174.640 1516.040 ;
        RECT 4.400 1509.920 1174.640 1511.320 ;
        RECT 4.000 1505.200 1174.640 1509.920 ;
        RECT 4.400 1503.800 1174.640 1505.200 ;
        RECT 4.000 1499.080 1174.640 1503.800 ;
        RECT 4.400 1497.680 1174.640 1499.080 ;
        RECT 4.000 1492.960 1174.640 1497.680 ;
        RECT 4.400 1491.560 1174.640 1492.960 ;
        RECT 4.000 1486.840 1174.640 1491.560 ;
        RECT 4.400 1485.440 1174.640 1486.840 ;
        RECT 4.000 1481.400 1174.640 1485.440 ;
        RECT 4.400 1480.000 1174.640 1481.400 ;
        RECT 4.000 1475.280 1174.640 1480.000 ;
        RECT 4.400 1473.880 1174.640 1475.280 ;
        RECT 4.000 1469.160 1174.640 1473.880 ;
        RECT 4.400 1467.760 1174.640 1469.160 ;
        RECT 4.000 1463.040 1174.640 1467.760 ;
        RECT 4.400 1461.640 1174.640 1463.040 ;
        RECT 4.000 1456.920 1174.640 1461.640 ;
        RECT 4.400 1455.520 1174.640 1456.920 ;
        RECT 4.000 1450.800 1174.640 1455.520 ;
        RECT 4.400 1449.400 1174.640 1450.800 ;
        RECT 4.000 1444.680 1174.640 1449.400 ;
        RECT 4.400 1443.280 1174.640 1444.680 ;
        RECT 4.000 1438.560 1174.640 1443.280 ;
        RECT 4.400 1437.160 1174.640 1438.560 ;
        RECT 4.000 1432.440 1174.640 1437.160 ;
        RECT 4.400 1431.040 1174.640 1432.440 ;
        RECT 4.000 1426.320 1174.640 1431.040 ;
        RECT 4.400 1424.920 1174.640 1426.320 ;
        RECT 4.000 1420.200 1174.640 1424.920 ;
        RECT 4.400 1418.800 1174.640 1420.200 ;
        RECT 4.000 1414.080 1174.640 1418.800 ;
        RECT 4.400 1412.680 1174.640 1414.080 ;
        RECT 4.000 1407.960 1174.640 1412.680 ;
        RECT 4.400 1406.560 1174.640 1407.960 ;
        RECT 4.000 1401.840 1174.640 1406.560 ;
        RECT 4.400 1400.440 1174.640 1401.840 ;
        RECT 4.000 1395.720 1174.640 1400.440 ;
        RECT 4.400 1394.320 1174.640 1395.720 ;
        RECT 4.000 1389.600 1174.640 1394.320 ;
        RECT 4.400 1388.200 1174.640 1389.600 ;
        RECT 4.000 1383.480 1174.640 1388.200 ;
        RECT 4.400 1382.080 1174.640 1383.480 ;
        RECT 4.000 1378.040 1174.640 1382.080 ;
        RECT 4.400 1376.640 1174.640 1378.040 ;
        RECT 4.000 1371.920 1174.640 1376.640 ;
        RECT 4.400 1370.520 1174.640 1371.920 ;
        RECT 4.000 1365.800 1174.640 1370.520 ;
        RECT 4.400 1364.400 1174.640 1365.800 ;
        RECT 4.000 1359.680 1174.640 1364.400 ;
        RECT 4.400 1358.280 1174.640 1359.680 ;
        RECT 4.000 1353.560 1174.640 1358.280 ;
        RECT 4.400 1352.160 1174.640 1353.560 ;
        RECT 4.000 1347.440 1174.640 1352.160 ;
        RECT 4.400 1346.040 1174.640 1347.440 ;
        RECT 4.000 1341.320 1174.640 1346.040 ;
        RECT 4.400 1339.920 1174.640 1341.320 ;
        RECT 4.000 1335.200 1174.640 1339.920 ;
        RECT 4.400 1333.800 1174.640 1335.200 ;
        RECT 4.000 1329.080 1174.640 1333.800 ;
        RECT 4.400 1327.680 1174.640 1329.080 ;
        RECT 4.000 1322.960 1174.640 1327.680 ;
        RECT 4.400 1321.560 1174.640 1322.960 ;
        RECT 4.000 1316.840 1174.640 1321.560 ;
        RECT 4.400 1315.440 1174.640 1316.840 ;
        RECT 4.000 1310.720 1174.640 1315.440 ;
        RECT 4.400 1309.320 1174.640 1310.720 ;
        RECT 4.000 1304.600 1174.640 1309.320 ;
        RECT 4.400 1303.200 1174.640 1304.600 ;
        RECT 4.000 1298.480 1174.640 1303.200 ;
        RECT 4.400 1297.080 1174.640 1298.480 ;
        RECT 4.000 1292.360 1174.640 1297.080 ;
        RECT 4.400 1290.960 1174.640 1292.360 ;
        RECT 4.000 1286.240 1174.640 1290.960 ;
        RECT 4.400 1284.840 1174.640 1286.240 ;
        RECT 4.000 1280.120 1174.640 1284.840 ;
        RECT 4.400 1278.720 1174.640 1280.120 ;
        RECT 4.000 1274.000 1174.640 1278.720 ;
        RECT 4.400 1272.600 1174.640 1274.000 ;
        RECT 4.000 1268.560 1174.640 1272.600 ;
        RECT 4.400 1267.160 1174.640 1268.560 ;
        RECT 4.000 1262.440 1174.640 1267.160 ;
        RECT 4.400 1261.040 1174.640 1262.440 ;
        RECT 4.000 1256.320 1174.640 1261.040 ;
        RECT 4.400 1254.920 1174.640 1256.320 ;
        RECT 4.000 1250.200 1174.640 1254.920 ;
        RECT 4.400 1248.800 1174.640 1250.200 ;
        RECT 4.000 1244.080 1174.640 1248.800 ;
        RECT 4.400 1242.680 1174.640 1244.080 ;
        RECT 4.000 1237.960 1174.640 1242.680 ;
        RECT 4.400 1236.560 1174.640 1237.960 ;
        RECT 4.000 1231.840 1174.640 1236.560 ;
        RECT 4.400 1230.440 1174.640 1231.840 ;
        RECT 4.000 1225.720 1174.640 1230.440 ;
        RECT 4.400 1224.320 1174.640 1225.720 ;
        RECT 4.000 1219.600 1174.640 1224.320 ;
        RECT 4.400 1218.200 1174.640 1219.600 ;
        RECT 4.000 1213.480 1174.640 1218.200 ;
        RECT 4.400 1212.080 1174.640 1213.480 ;
        RECT 4.000 1207.360 1174.640 1212.080 ;
        RECT 4.400 1205.960 1174.640 1207.360 ;
        RECT 4.000 1201.240 1174.640 1205.960 ;
        RECT 4.400 1199.840 1174.640 1201.240 ;
        RECT 4.000 1195.120 1174.640 1199.840 ;
        RECT 4.400 1193.720 1174.640 1195.120 ;
        RECT 4.000 1189.000 1174.640 1193.720 ;
        RECT 4.400 1187.600 1174.640 1189.000 ;
        RECT 4.000 1182.880 1174.640 1187.600 ;
        RECT 4.400 1181.480 1174.640 1182.880 ;
        RECT 4.000 1176.760 1174.640 1181.480 ;
        RECT 4.400 1175.360 1174.640 1176.760 ;
        RECT 4.000 1170.640 1174.640 1175.360 ;
        RECT 4.400 1169.240 1174.640 1170.640 ;
        RECT 4.000 1165.200 1174.640 1169.240 ;
        RECT 4.400 1163.800 1174.640 1165.200 ;
        RECT 4.000 1159.080 1174.640 1163.800 ;
        RECT 4.400 1157.680 1174.640 1159.080 ;
        RECT 4.000 1152.960 1174.640 1157.680 ;
        RECT 4.400 1151.560 1174.640 1152.960 ;
        RECT 4.000 1146.840 1174.640 1151.560 ;
        RECT 4.400 1145.440 1174.640 1146.840 ;
        RECT 4.000 1140.720 1174.640 1145.440 ;
        RECT 4.400 1139.320 1174.640 1140.720 ;
        RECT 4.000 1134.600 1174.640 1139.320 ;
        RECT 4.400 1133.200 1174.640 1134.600 ;
        RECT 4.000 1128.480 1174.640 1133.200 ;
        RECT 4.400 1127.080 1174.640 1128.480 ;
        RECT 4.000 1122.360 1174.640 1127.080 ;
        RECT 4.400 1120.960 1174.640 1122.360 ;
        RECT 4.000 1116.240 1174.640 1120.960 ;
        RECT 4.400 1114.840 1174.640 1116.240 ;
        RECT 4.000 1110.120 1174.640 1114.840 ;
        RECT 4.400 1108.720 1174.640 1110.120 ;
        RECT 4.000 1104.000 1174.640 1108.720 ;
        RECT 4.400 1102.600 1174.640 1104.000 ;
        RECT 4.000 1097.880 1174.640 1102.600 ;
        RECT 4.400 1096.480 1174.640 1097.880 ;
        RECT 4.000 1091.760 1174.640 1096.480 ;
        RECT 4.400 1090.360 1174.640 1091.760 ;
        RECT 4.000 1085.640 1174.640 1090.360 ;
        RECT 4.400 1084.240 1174.640 1085.640 ;
        RECT 4.000 1079.520 1174.640 1084.240 ;
        RECT 4.400 1078.120 1174.640 1079.520 ;
        RECT 4.000 1073.400 1174.640 1078.120 ;
        RECT 4.400 1072.000 1174.640 1073.400 ;
        RECT 4.000 1067.280 1174.640 1072.000 ;
        RECT 4.400 1065.880 1174.640 1067.280 ;
        RECT 4.000 1061.840 1174.640 1065.880 ;
        RECT 4.400 1060.440 1174.640 1061.840 ;
        RECT 4.000 1055.720 1174.640 1060.440 ;
        RECT 4.400 1054.320 1174.640 1055.720 ;
        RECT 4.000 1049.600 1174.640 1054.320 ;
        RECT 4.400 1048.200 1174.640 1049.600 ;
        RECT 4.000 1043.480 1174.640 1048.200 ;
        RECT 4.400 1042.080 1174.640 1043.480 ;
        RECT 4.000 1037.360 1174.640 1042.080 ;
        RECT 4.400 1035.960 1174.640 1037.360 ;
        RECT 4.000 1031.240 1174.640 1035.960 ;
        RECT 4.400 1029.840 1174.640 1031.240 ;
        RECT 4.000 1025.120 1174.640 1029.840 ;
        RECT 4.400 1023.720 1174.640 1025.120 ;
        RECT 4.000 1019.000 1174.640 1023.720 ;
        RECT 4.400 1017.600 1174.640 1019.000 ;
        RECT 4.000 1012.880 1174.640 1017.600 ;
        RECT 4.400 1011.480 1174.640 1012.880 ;
        RECT 4.000 1006.760 1174.640 1011.480 ;
        RECT 4.400 1005.360 1174.640 1006.760 ;
        RECT 4.000 1000.640 1174.640 1005.360 ;
        RECT 4.400 999.240 1174.640 1000.640 ;
        RECT 4.000 994.520 1174.640 999.240 ;
        RECT 4.400 993.120 1174.640 994.520 ;
        RECT 4.000 988.400 1174.640 993.120 ;
        RECT 4.400 987.000 1174.640 988.400 ;
        RECT 4.000 982.280 1174.640 987.000 ;
        RECT 4.400 980.880 1174.640 982.280 ;
        RECT 4.000 976.160 1174.640 980.880 ;
        RECT 4.400 974.760 1174.640 976.160 ;
        RECT 4.000 970.040 1174.640 974.760 ;
        RECT 4.400 968.640 1174.640 970.040 ;
        RECT 4.000 963.920 1174.640 968.640 ;
        RECT 4.400 962.520 1174.640 963.920 ;
        RECT 4.000 957.800 1174.640 962.520 ;
        RECT 4.400 956.400 1174.640 957.800 ;
        RECT 4.000 952.360 1174.640 956.400 ;
        RECT 4.400 950.960 1174.640 952.360 ;
        RECT 4.000 946.240 1174.640 950.960 ;
        RECT 4.400 944.840 1174.640 946.240 ;
        RECT 4.000 940.120 1174.640 944.840 ;
        RECT 4.400 938.720 1174.640 940.120 ;
        RECT 4.000 934.000 1174.640 938.720 ;
        RECT 4.400 932.600 1174.640 934.000 ;
        RECT 4.000 927.880 1174.640 932.600 ;
        RECT 4.400 926.480 1174.640 927.880 ;
        RECT 4.000 921.760 1174.640 926.480 ;
        RECT 4.400 920.360 1174.640 921.760 ;
        RECT 4.000 915.640 1174.640 920.360 ;
        RECT 4.400 914.240 1174.640 915.640 ;
        RECT 4.000 909.520 1174.640 914.240 ;
        RECT 4.400 908.120 1174.640 909.520 ;
        RECT 4.000 903.400 1174.640 908.120 ;
        RECT 4.400 902.000 1174.640 903.400 ;
        RECT 4.000 897.280 1174.640 902.000 ;
        RECT 4.400 895.880 1174.640 897.280 ;
        RECT 4.000 891.160 1174.640 895.880 ;
        RECT 4.400 889.760 1174.640 891.160 ;
        RECT 4.000 885.040 1174.640 889.760 ;
        RECT 4.400 883.640 1174.640 885.040 ;
        RECT 4.000 878.920 1174.640 883.640 ;
        RECT 4.400 877.520 1174.640 878.920 ;
        RECT 4.000 872.800 1174.640 877.520 ;
        RECT 4.400 871.400 1174.640 872.800 ;
        RECT 4.000 866.680 1174.640 871.400 ;
        RECT 4.400 865.280 1174.640 866.680 ;
        RECT 4.000 860.560 1174.640 865.280 ;
        RECT 4.400 859.160 1174.640 860.560 ;
        RECT 4.000 854.440 1174.640 859.160 ;
        RECT 4.400 853.040 1174.640 854.440 ;
        RECT 4.000 849.000 1174.640 853.040 ;
        RECT 4.400 847.600 1174.640 849.000 ;
        RECT 4.000 842.880 1174.640 847.600 ;
        RECT 4.400 841.480 1174.640 842.880 ;
        RECT 4.000 836.760 1174.640 841.480 ;
        RECT 4.400 835.360 1174.640 836.760 ;
        RECT 4.000 830.640 1174.640 835.360 ;
        RECT 4.400 829.240 1174.640 830.640 ;
        RECT 4.000 824.520 1174.640 829.240 ;
        RECT 4.400 823.120 1174.640 824.520 ;
        RECT 4.000 818.400 1174.640 823.120 ;
        RECT 4.400 817.000 1174.640 818.400 ;
        RECT 4.000 812.280 1174.640 817.000 ;
        RECT 4.400 810.880 1174.640 812.280 ;
        RECT 4.000 806.160 1174.640 810.880 ;
        RECT 4.400 804.760 1174.640 806.160 ;
        RECT 4.000 800.040 1174.640 804.760 ;
        RECT 4.400 798.640 1174.640 800.040 ;
        RECT 4.000 793.920 1174.640 798.640 ;
        RECT 4.400 792.520 1174.640 793.920 ;
        RECT 4.000 787.800 1174.640 792.520 ;
        RECT 4.400 786.400 1174.640 787.800 ;
        RECT 4.000 781.680 1174.640 786.400 ;
        RECT 4.400 780.280 1174.640 781.680 ;
        RECT 4.000 775.560 1174.640 780.280 ;
        RECT 4.400 774.160 1174.640 775.560 ;
        RECT 4.000 769.440 1174.640 774.160 ;
        RECT 4.400 768.040 1174.640 769.440 ;
        RECT 4.000 763.320 1174.640 768.040 ;
        RECT 4.400 761.920 1174.640 763.320 ;
        RECT 4.000 757.200 1174.640 761.920 ;
        RECT 4.400 755.800 1174.640 757.200 ;
        RECT 4.000 751.080 1174.640 755.800 ;
        RECT 4.400 749.680 1174.640 751.080 ;
        RECT 4.000 744.960 1174.640 749.680 ;
        RECT 4.400 743.560 1174.640 744.960 ;
        RECT 4.000 739.520 1174.640 743.560 ;
        RECT 4.400 738.120 1174.640 739.520 ;
        RECT 4.000 733.400 1174.640 738.120 ;
        RECT 4.400 732.000 1174.640 733.400 ;
        RECT 4.000 727.280 1174.640 732.000 ;
        RECT 4.400 725.880 1174.640 727.280 ;
        RECT 4.000 721.160 1174.640 725.880 ;
        RECT 4.400 719.760 1174.640 721.160 ;
        RECT 4.000 715.040 1174.640 719.760 ;
        RECT 4.400 713.640 1174.640 715.040 ;
        RECT 4.000 708.920 1174.640 713.640 ;
        RECT 4.400 707.520 1174.640 708.920 ;
        RECT 4.000 702.800 1174.640 707.520 ;
        RECT 4.400 701.400 1174.640 702.800 ;
        RECT 4.000 696.680 1174.640 701.400 ;
        RECT 4.400 695.280 1174.640 696.680 ;
        RECT 4.000 690.560 1174.640 695.280 ;
        RECT 4.400 689.160 1174.640 690.560 ;
        RECT 4.000 684.440 1174.640 689.160 ;
        RECT 4.400 683.040 1174.640 684.440 ;
        RECT 4.000 678.320 1174.640 683.040 ;
        RECT 4.400 676.920 1174.640 678.320 ;
        RECT 4.000 672.200 1174.640 676.920 ;
        RECT 4.400 670.800 1174.640 672.200 ;
        RECT 4.000 666.080 1174.640 670.800 ;
        RECT 4.400 664.680 1174.640 666.080 ;
        RECT 4.000 659.960 1174.640 664.680 ;
        RECT 4.400 658.560 1174.640 659.960 ;
        RECT 4.000 653.840 1174.640 658.560 ;
        RECT 4.400 652.440 1174.640 653.840 ;
        RECT 4.000 647.720 1174.640 652.440 ;
        RECT 4.400 646.320 1174.640 647.720 ;
        RECT 4.000 641.600 1174.640 646.320 ;
        RECT 4.400 640.200 1174.640 641.600 ;
        RECT 4.000 636.160 1174.640 640.200 ;
        RECT 4.400 634.760 1174.640 636.160 ;
        RECT 4.000 630.040 1174.640 634.760 ;
        RECT 4.400 628.640 1174.640 630.040 ;
        RECT 4.000 623.920 1174.640 628.640 ;
        RECT 4.400 622.520 1174.640 623.920 ;
        RECT 4.000 617.800 1174.640 622.520 ;
        RECT 4.400 616.400 1174.640 617.800 ;
        RECT 4.000 611.680 1174.640 616.400 ;
        RECT 4.400 610.280 1174.640 611.680 ;
        RECT 4.000 605.560 1174.640 610.280 ;
        RECT 4.400 604.160 1174.640 605.560 ;
        RECT 4.000 599.440 1174.640 604.160 ;
        RECT 4.400 598.040 1174.640 599.440 ;
        RECT 4.000 593.320 1174.640 598.040 ;
        RECT 4.400 591.920 1174.640 593.320 ;
        RECT 4.000 587.200 1174.640 591.920 ;
        RECT 4.400 585.800 1174.640 587.200 ;
        RECT 4.000 581.080 1174.640 585.800 ;
        RECT 4.400 579.680 1174.640 581.080 ;
        RECT 4.000 574.960 1174.640 579.680 ;
        RECT 4.400 573.560 1174.640 574.960 ;
        RECT 4.000 568.840 1174.640 573.560 ;
        RECT 4.400 567.440 1174.640 568.840 ;
        RECT 4.000 562.720 1174.640 567.440 ;
        RECT 4.400 561.320 1174.640 562.720 ;
        RECT 4.000 556.600 1174.640 561.320 ;
        RECT 4.400 555.200 1174.640 556.600 ;
        RECT 4.000 550.480 1174.640 555.200 ;
        RECT 4.400 549.080 1174.640 550.480 ;
        RECT 4.000 544.360 1174.640 549.080 ;
        RECT 4.400 542.960 1174.640 544.360 ;
        RECT 4.000 538.240 1174.640 542.960 ;
        RECT 4.400 536.840 1174.640 538.240 ;
        RECT 4.000 532.800 1174.640 536.840 ;
        RECT 4.400 531.400 1174.640 532.800 ;
        RECT 4.000 526.680 1174.640 531.400 ;
        RECT 4.400 525.280 1174.640 526.680 ;
        RECT 4.000 520.560 1174.640 525.280 ;
        RECT 4.400 519.160 1174.640 520.560 ;
        RECT 4.000 514.440 1174.640 519.160 ;
        RECT 4.400 513.040 1174.640 514.440 ;
        RECT 4.000 508.320 1174.640 513.040 ;
        RECT 4.400 506.920 1174.640 508.320 ;
        RECT 4.000 502.200 1174.640 506.920 ;
        RECT 4.400 500.800 1174.640 502.200 ;
        RECT 4.000 496.080 1174.640 500.800 ;
        RECT 4.400 494.680 1174.640 496.080 ;
        RECT 4.000 489.960 1174.640 494.680 ;
        RECT 4.400 488.560 1174.640 489.960 ;
        RECT 4.000 483.840 1174.640 488.560 ;
        RECT 4.400 482.440 1174.640 483.840 ;
        RECT 4.000 477.720 1174.640 482.440 ;
        RECT 4.400 476.320 1174.640 477.720 ;
        RECT 4.000 471.600 1174.640 476.320 ;
        RECT 4.400 470.200 1174.640 471.600 ;
        RECT 4.000 465.480 1174.640 470.200 ;
        RECT 4.400 464.080 1174.640 465.480 ;
        RECT 4.000 459.360 1174.640 464.080 ;
        RECT 4.400 457.960 1174.640 459.360 ;
        RECT 4.000 453.240 1174.640 457.960 ;
        RECT 4.400 451.840 1174.640 453.240 ;
        RECT 4.000 447.120 1174.640 451.840 ;
        RECT 4.400 445.720 1174.640 447.120 ;
        RECT 4.000 441.000 1174.640 445.720 ;
        RECT 4.400 439.600 1174.640 441.000 ;
        RECT 4.000 434.880 1174.640 439.600 ;
        RECT 4.400 433.480 1174.640 434.880 ;
        RECT 4.000 428.760 1174.640 433.480 ;
        RECT 4.400 427.360 1174.640 428.760 ;
        RECT 4.000 423.320 1174.640 427.360 ;
        RECT 4.400 421.920 1174.640 423.320 ;
        RECT 4.000 417.200 1174.640 421.920 ;
        RECT 4.400 415.800 1174.640 417.200 ;
        RECT 4.000 411.080 1174.640 415.800 ;
        RECT 4.400 409.680 1174.640 411.080 ;
        RECT 4.000 404.960 1174.640 409.680 ;
        RECT 4.400 403.560 1174.640 404.960 ;
        RECT 4.000 398.840 1174.640 403.560 ;
        RECT 4.400 397.440 1174.640 398.840 ;
        RECT 4.000 392.720 1174.640 397.440 ;
        RECT 4.400 391.320 1174.640 392.720 ;
        RECT 4.000 386.600 1174.640 391.320 ;
        RECT 4.400 385.200 1174.640 386.600 ;
        RECT 4.000 380.480 1174.640 385.200 ;
        RECT 4.400 379.080 1174.640 380.480 ;
        RECT 4.000 374.360 1174.640 379.080 ;
        RECT 4.400 372.960 1174.640 374.360 ;
        RECT 4.000 368.240 1174.640 372.960 ;
        RECT 4.400 366.840 1174.640 368.240 ;
        RECT 4.000 362.120 1174.640 366.840 ;
        RECT 4.400 360.720 1174.640 362.120 ;
        RECT 4.000 356.000 1174.640 360.720 ;
        RECT 4.400 354.600 1174.640 356.000 ;
        RECT 4.000 349.880 1174.640 354.600 ;
        RECT 4.400 348.480 1174.640 349.880 ;
        RECT 4.000 343.760 1174.640 348.480 ;
        RECT 4.400 342.360 1174.640 343.760 ;
        RECT 4.000 337.640 1174.640 342.360 ;
        RECT 4.400 336.240 1174.640 337.640 ;
        RECT 4.000 331.520 1174.640 336.240 ;
        RECT 4.400 330.120 1174.640 331.520 ;
        RECT 4.000 325.400 1174.640 330.120 ;
        RECT 4.400 324.000 1174.640 325.400 ;
        RECT 4.000 319.960 1174.640 324.000 ;
        RECT 4.400 318.560 1174.640 319.960 ;
        RECT 4.000 313.840 1174.640 318.560 ;
        RECT 4.400 312.440 1174.640 313.840 ;
        RECT 4.000 307.720 1174.640 312.440 ;
        RECT 4.400 306.320 1174.640 307.720 ;
        RECT 4.000 301.600 1174.640 306.320 ;
        RECT 4.400 300.200 1174.640 301.600 ;
        RECT 4.000 295.480 1174.640 300.200 ;
        RECT 4.400 294.080 1174.640 295.480 ;
        RECT 4.000 289.360 1174.640 294.080 ;
        RECT 4.400 287.960 1174.640 289.360 ;
        RECT 4.000 283.240 1174.640 287.960 ;
        RECT 4.400 281.840 1174.640 283.240 ;
        RECT 4.000 277.120 1174.640 281.840 ;
        RECT 4.400 275.720 1174.640 277.120 ;
        RECT 4.000 271.000 1174.640 275.720 ;
        RECT 4.400 269.600 1174.640 271.000 ;
        RECT 4.000 264.880 1174.640 269.600 ;
        RECT 4.400 263.480 1174.640 264.880 ;
        RECT 4.000 258.760 1174.640 263.480 ;
        RECT 4.400 257.360 1174.640 258.760 ;
        RECT 4.000 252.640 1174.640 257.360 ;
        RECT 4.400 251.240 1174.640 252.640 ;
        RECT 4.000 246.520 1174.640 251.240 ;
        RECT 4.400 245.120 1174.640 246.520 ;
        RECT 4.000 240.400 1174.640 245.120 ;
        RECT 4.400 239.000 1174.640 240.400 ;
        RECT 4.000 234.280 1174.640 239.000 ;
        RECT 4.400 232.880 1174.640 234.280 ;
        RECT 4.000 228.160 1174.640 232.880 ;
        RECT 4.400 226.760 1174.640 228.160 ;
        RECT 4.000 222.040 1174.640 226.760 ;
        RECT 4.400 220.640 1174.640 222.040 ;
        RECT 4.000 215.920 1174.640 220.640 ;
        RECT 4.400 214.520 1174.640 215.920 ;
        RECT 4.000 210.480 1174.640 214.520 ;
        RECT 4.400 209.080 1174.640 210.480 ;
        RECT 4.000 204.360 1174.640 209.080 ;
        RECT 4.400 202.960 1174.640 204.360 ;
        RECT 4.000 198.240 1174.640 202.960 ;
        RECT 4.400 196.840 1174.640 198.240 ;
        RECT 4.000 192.120 1174.640 196.840 ;
        RECT 4.400 190.720 1174.640 192.120 ;
        RECT 4.000 186.000 1174.640 190.720 ;
        RECT 4.400 184.600 1174.640 186.000 ;
        RECT 4.000 179.880 1174.640 184.600 ;
        RECT 4.400 178.480 1174.640 179.880 ;
        RECT 4.000 173.760 1174.640 178.480 ;
        RECT 4.400 172.360 1174.640 173.760 ;
        RECT 4.000 167.640 1174.640 172.360 ;
        RECT 4.400 166.240 1174.640 167.640 ;
        RECT 4.000 161.520 1174.640 166.240 ;
        RECT 4.400 160.120 1174.640 161.520 ;
        RECT 4.000 155.400 1174.640 160.120 ;
        RECT 4.400 154.000 1174.640 155.400 ;
        RECT 4.000 149.280 1174.640 154.000 ;
        RECT 4.400 147.880 1174.640 149.280 ;
        RECT 4.000 143.160 1174.640 147.880 ;
        RECT 4.400 141.760 1174.640 143.160 ;
        RECT 4.000 137.040 1174.640 141.760 ;
        RECT 4.400 135.640 1174.640 137.040 ;
        RECT 4.000 130.920 1174.640 135.640 ;
        RECT 4.400 129.520 1174.640 130.920 ;
        RECT 4.000 124.800 1174.640 129.520 ;
        RECT 4.400 123.400 1174.640 124.800 ;
        RECT 4.000 118.680 1174.640 123.400 ;
        RECT 4.400 117.280 1174.640 118.680 ;
        RECT 4.000 112.560 1174.640 117.280 ;
        RECT 4.400 111.160 1174.640 112.560 ;
        RECT 4.000 107.120 1174.640 111.160 ;
        RECT 4.400 105.720 1174.640 107.120 ;
        RECT 4.000 101.000 1174.640 105.720 ;
        RECT 4.400 99.600 1174.640 101.000 ;
        RECT 4.000 94.880 1174.640 99.600 ;
        RECT 4.400 93.480 1174.640 94.880 ;
        RECT 4.000 88.760 1174.640 93.480 ;
        RECT 4.400 87.360 1174.640 88.760 ;
        RECT 4.000 82.640 1174.640 87.360 ;
        RECT 4.400 81.240 1174.640 82.640 ;
        RECT 4.000 76.520 1174.640 81.240 ;
        RECT 4.400 75.120 1174.640 76.520 ;
        RECT 4.000 70.400 1174.640 75.120 ;
        RECT 4.400 69.000 1174.640 70.400 ;
        RECT 4.000 64.280 1174.640 69.000 ;
        RECT 4.400 62.880 1174.640 64.280 ;
        RECT 4.000 58.160 1174.640 62.880 ;
        RECT 4.400 56.760 1174.640 58.160 ;
        RECT 4.000 52.040 1174.640 56.760 ;
        RECT 4.400 50.640 1174.640 52.040 ;
        RECT 4.000 45.920 1174.640 50.640 ;
        RECT 4.400 44.520 1174.640 45.920 ;
        RECT 4.000 39.800 1174.640 44.520 ;
        RECT 4.400 38.400 1174.640 39.800 ;
        RECT 4.000 33.680 1174.640 38.400 ;
        RECT 4.400 32.280 1174.640 33.680 ;
        RECT 4.000 27.560 1174.640 32.280 ;
        RECT 4.400 26.160 1174.640 27.560 ;
        RECT 4.000 21.440 1174.640 26.160 ;
        RECT 4.400 20.040 1174.640 21.440 ;
        RECT 4.000 15.320 1174.640 20.040 ;
        RECT 4.400 13.920 1174.640 15.320 ;
        RECT 4.000 9.200 1174.640 13.920 ;
        RECT 4.400 7.800 1174.640 9.200 ;
        RECT 4.000 3.760 1174.640 7.800 ;
        RECT 4.400 2.895 1174.640 3.760 ;
      LAYER met4 ;
        RECT 7.655 11.735 20.640 1754.905 ;
        RECT 23.040 11.735 97.440 1754.905 ;
        RECT 99.840 11.735 174.240 1754.905 ;
        RECT 176.640 11.735 251.040 1754.905 ;
        RECT 253.440 11.735 327.840 1754.905 ;
        RECT 330.240 11.735 404.640 1754.905 ;
        RECT 407.040 11.735 481.440 1754.905 ;
        RECT 483.840 11.735 558.240 1754.905 ;
        RECT 560.640 11.735 635.040 1754.905 ;
        RECT 637.440 11.735 711.840 1754.905 ;
        RECT 714.240 11.735 788.640 1754.905 ;
        RECT 791.040 11.735 817.585 1754.905 ;
  END
END c0_system
END LIBRARY


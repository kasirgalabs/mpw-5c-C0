VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO c0_system
  CLASS BLOCK ;
  FOREIGN c0_system ;
  ORIGIN 0.000 0.000 ;
  SIZE 1600.000 BY 1600.000 ;
  PIN bb_addr0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 715.400 4.000 716.000 ;
    END
  END bb_addr0[0]
  PIN bb_addr0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1007.120 4.000 1007.720 ;
    END
  END bb_addr0[10]
  PIN bb_addr0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1034.320 4.000 1034.920 ;
    END
  END bb_addr0[11]
  PIN bb_addr0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1061.520 4.000 1062.120 ;
    END
  END bb_addr0[12]
  PIN bb_addr0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1088.040 4.000 1088.640 ;
    END
  END bb_addr0[13]
  PIN bb_addr0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1115.240 4.000 1115.840 ;
    END
  END bb_addr0[14]
  PIN bb_addr0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1142.440 4.000 1143.040 ;
    END
  END bb_addr0[15]
  PIN bb_addr0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1169.640 4.000 1170.240 ;
    END
  END bb_addr0[16]
  PIN bb_addr0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1196.160 4.000 1196.760 ;
    END
  END bb_addr0[17]
  PIN bb_addr0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1223.360 4.000 1223.960 ;
    END
  END bb_addr0[18]
  PIN bb_addr0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1250.560 4.000 1251.160 ;
    END
  END bb_addr0[19]
  PIN bb_addr0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 748.040 4.000 748.640 ;
    END
  END bb_addr0[1]
  PIN bb_addr0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1277.760 4.000 1278.360 ;
    END
  END bb_addr0[20]
  PIN bb_addr0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1304.280 4.000 1304.880 ;
    END
  END bb_addr0[21]
  PIN bb_addr0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1331.480 4.000 1332.080 ;
    END
  END bb_addr0[22]
  PIN bb_addr0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1358.680 4.000 1359.280 ;
    END
  END bb_addr0[23]
  PIN bb_addr0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1385.880 4.000 1386.480 ;
    END
  END bb_addr0[24]
  PIN bb_addr0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1412.400 4.000 1413.000 ;
    END
  END bb_addr0[25]
  PIN bb_addr0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1439.600 4.000 1440.200 ;
    END
  END bb_addr0[26]
  PIN bb_addr0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1466.800 4.000 1467.400 ;
    END
  END bb_addr0[27]
  PIN bb_addr0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1494.000 4.000 1494.600 ;
    END
  END bb_addr0[28]
  PIN bb_addr0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1520.520 4.000 1521.120 ;
    END
  END bb_addr0[29]
  PIN bb_addr0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 780.000 4.000 780.600 ;
    END
  END bb_addr0[2]
  PIN bb_addr0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1547.720 4.000 1548.320 ;
    END
  END bb_addr0[30]
  PIN bb_addr0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1574.920 4.000 1575.520 ;
    END
  END bb_addr0[31]
  PIN bb_addr0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 812.640 4.000 813.240 ;
    END
  END bb_addr0[3]
  PIN bb_addr0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 845.280 4.000 845.880 ;
    END
  END bb_addr0[4]
  PIN bb_addr0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 871.800 4.000 872.400 ;
    END
  END bb_addr0[5]
  PIN bb_addr0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 899.000 4.000 899.600 ;
    END
  END bb_addr0[6]
  PIN bb_addr0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 926.200 4.000 926.800 ;
    END
  END bb_addr0[7]
  PIN bb_addr0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 953.400 4.000 954.000 ;
    END
  END bb_addr0[8]
  PIN bb_addr0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 979.920 4.000 980.520 ;
    END
  END bb_addr0[9]
  PIN bb_addr1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 720.840 4.000 721.440 ;
    END
  END bb_addr1[0]
  PIN bb_addr1[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1012.560 4.000 1013.160 ;
    END
  END bb_addr1[10]
  PIN bb_addr1[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1039.760 4.000 1040.360 ;
    END
  END bb_addr1[11]
  PIN bb_addr1[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1066.960 4.000 1067.560 ;
    END
  END bb_addr1[12]
  PIN bb_addr1[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1093.480 4.000 1094.080 ;
    END
  END bb_addr1[13]
  PIN bb_addr1[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1120.680 4.000 1121.280 ;
    END
  END bb_addr1[14]
  PIN bb_addr1[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1147.880 4.000 1148.480 ;
    END
  END bb_addr1[15]
  PIN bb_addr1[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1175.080 4.000 1175.680 ;
    END
  END bb_addr1[16]
  PIN bb_addr1[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1201.600 4.000 1202.200 ;
    END
  END bb_addr1[17]
  PIN bb_addr1[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1228.800 4.000 1229.400 ;
    END
  END bb_addr1[18]
  PIN bb_addr1[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1256.000 4.000 1256.600 ;
    END
  END bb_addr1[19]
  PIN bb_addr1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 752.800 4.000 753.400 ;
    END
  END bb_addr1[1]
  PIN bb_addr1[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1282.520 4.000 1283.120 ;
    END
  END bb_addr1[20]
  PIN bb_addr1[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1309.720 4.000 1310.320 ;
    END
  END bb_addr1[21]
  PIN bb_addr1[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1336.920 4.000 1337.520 ;
    END
  END bb_addr1[22]
  PIN bb_addr1[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1364.120 4.000 1364.720 ;
    END
  END bb_addr1[23]
  PIN bb_addr1[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1390.640 4.000 1391.240 ;
    END
  END bb_addr1[24]
  PIN bb_addr1[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1417.840 4.000 1418.440 ;
    END
  END bb_addr1[25]
  PIN bb_addr1[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1445.040 4.000 1445.640 ;
    END
  END bb_addr1[26]
  PIN bb_addr1[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1472.240 4.000 1472.840 ;
    END
  END bb_addr1[27]
  PIN bb_addr1[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1498.760 4.000 1499.360 ;
    END
  END bb_addr1[28]
  PIN bb_addr1[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1525.960 4.000 1526.560 ;
    END
  END bb_addr1[29]
  PIN bb_addr1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 785.440 4.000 786.040 ;
    END
  END bb_addr1[2]
  PIN bb_addr1[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1553.160 4.000 1553.760 ;
    END
  END bb_addr1[30]
  PIN bb_addr1[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1580.360 4.000 1580.960 ;
    END
  END bb_addr1[31]
  PIN bb_addr1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 818.080 4.000 818.680 ;
    END
  END bb_addr1[3]
  PIN bb_addr1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 850.720 4.000 851.320 ;
    END
  END bb_addr1[4]
  PIN bb_addr1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 877.240 4.000 877.840 ;
    END
  END bb_addr1[5]
  PIN bb_addr1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 904.440 4.000 905.040 ;
    END
  END bb_addr1[6]
  PIN bb_addr1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 931.640 4.000 932.240 ;
    END
  END bb_addr1[7]
  PIN bb_addr1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 958.840 4.000 959.440 ;
    END
  END bb_addr1[8]
  PIN bb_addr1[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 985.360 4.000 985.960 ;
    END
  END bb_addr1[9]
  PIN bb_csb0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 699.080 4.000 699.680 ;
    END
  END bb_csb0
  PIN bb_csb1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 704.520 4.000 705.120 ;
    END
  END bb_csb1
  PIN bb_din0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 726.280 4.000 726.880 ;
    END
  END bb_din0[0]
  PIN bb_din0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1018.000 4.000 1018.600 ;
    END
  END bb_din0[10]
  PIN bb_din0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1045.200 4.000 1045.800 ;
    END
  END bb_din0[11]
  PIN bb_din0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1071.720 4.000 1072.320 ;
    END
  END bb_din0[12]
  PIN bb_din0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1098.920 4.000 1099.520 ;
    END
  END bb_din0[13]
  PIN bb_din0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1126.120 4.000 1126.720 ;
    END
  END bb_din0[14]
  PIN bb_din0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1153.320 4.000 1153.920 ;
    END
  END bb_din0[15]
  PIN bb_din0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1179.840 4.000 1180.440 ;
    END
  END bb_din0[16]
  PIN bb_din0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1207.040 4.000 1207.640 ;
    END
  END bb_din0[17]
  PIN bb_din0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1234.240 4.000 1234.840 ;
    END
  END bb_din0[18]
  PIN bb_din0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1261.440 4.000 1262.040 ;
    END
  END bb_din0[19]
  PIN bb_din0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 758.240 4.000 758.840 ;
    END
  END bb_din0[1]
  PIN bb_din0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1287.960 4.000 1288.560 ;
    END
  END bb_din0[20]
  PIN bb_din0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1315.160 4.000 1315.760 ;
    END
  END bb_din0[21]
  PIN bb_din0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1342.360 4.000 1342.960 ;
    END
  END bb_din0[22]
  PIN bb_din0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1369.560 4.000 1370.160 ;
    END
  END bb_din0[23]
  PIN bb_din0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1396.080 4.000 1396.680 ;
    END
  END bb_din0[24]
  PIN bb_din0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1423.280 4.000 1423.880 ;
    END
  END bb_din0[25]
  PIN bb_din0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1450.480 4.000 1451.080 ;
    END
  END bb_din0[26]
  PIN bb_din0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1477.680 4.000 1478.280 ;
    END
  END bb_din0[27]
  PIN bb_din0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1504.200 4.000 1504.800 ;
    END
  END bb_din0[28]
  PIN bb_din0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1531.400 4.000 1532.000 ;
    END
  END bb_din0[29]
  PIN bb_din0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 790.880 4.000 791.480 ;
    END
  END bb_din0[2]
  PIN bb_din0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1558.600 4.000 1559.200 ;
    END
  END bb_din0[30]
  PIN bb_din0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1585.800 4.000 1586.400 ;
    END
  END bb_din0[31]
  PIN bb_din0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 823.520 4.000 824.120 ;
    END
  END bb_din0[3]
  PIN bb_din0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 855.480 4.000 856.080 ;
    END
  END bb_din0[4]
  PIN bb_din0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 882.680 4.000 883.280 ;
    END
  END bb_din0[5]
  PIN bb_din0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 909.880 4.000 910.480 ;
    END
  END bb_din0[6]
  PIN bb_din0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 937.080 4.000 937.680 ;
    END
  END bb_din0[7]
  PIN bb_din0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 963.600 4.000 964.200 ;
    END
  END bb_din0[8]
  PIN bb_din0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 990.800 4.000 991.400 ;
    END
  END bb_din0[9]
  PIN bb_dout0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 731.720 4.000 732.320 ;
    END
  END bb_dout0[0]
  PIN bb_dout0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1023.440 4.000 1024.040 ;
    END
  END bb_dout0[10]
  PIN bb_dout0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1050.640 4.000 1051.240 ;
    END
  END bb_dout0[11]
  PIN bb_dout0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1077.160 4.000 1077.760 ;
    END
  END bb_dout0[12]
  PIN bb_dout0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1104.360 4.000 1104.960 ;
    END
  END bb_dout0[13]
  PIN bb_dout0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1131.560 4.000 1132.160 ;
    END
  END bb_dout0[14]
  PIN bb_dout0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1158.760 4.000 1159.360 ;
    END
  END bb_dout0[15]
  PIN bb_dout0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1185.280 4.000 1185.880 ;
    END
  END bb_dout0[16]
  PIN bb_dout0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1212.480 4.000 1213.080 ;
    END
  END bb_dout0[17]
  PIN bb_dout0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1239.680 4.000 1240.280 ;
    END
  END bb_dout0[18]
  PIN bb_dout0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1266.880 4.000 1267.480 ;
    END
  END bb_dout0[19]
  PIN bb_dout0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 763.680 4.000 764.280 ;
    END
  END bb_dout0[1]
  PIN bb_dout0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1293.400 4.000 1294.000 ;
    END
  END bb_dout0[20]
  PIN bb_dout0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1320.600 4.000 1321.200 ;
    END
  END bb_dout0[21]
  PIN bb_dout0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1347.800 4.000 1348.400 ;
    END
  END bb_dout0[22]
  PIN bb_dout0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1375.000 4.000 1375.600 ;
    END
  END bb_dout0[23]
  PIN bb_dout0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1401.520 4.000 1402.120 ;
    END
  END bb_dout0[24]
  PIN bb_dout0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1428.720 4.000 1429.320 ;
    END
  END bb_dout0[25]
  PIN bb_dout0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1455.920 4.000 1456.520 ;
    END
  END bb_dout0[26]
  PIN bb_dout0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1483.120 4.000 1483.720 ;
    END
  END bb_dout0[27]
  PIN bb_dout0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1509.640 4.000 1510.240 ;
    END
  END bb_dout0[28]
  PIN bb_dout0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1536.840 4.000 1537.440 ;
    END
  END bb_dout0[29]
  PIN bb_dout0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 796.320 4.000 796.920 ;
    END
  END bb_dout0[2]
  PIN bb_dout0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1564.040 4.000 1564.640 ;
    END
  END bb_dout0[30]
  PIN bb_dout0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1591.240 4.000 1591.840 ;
    END
  END bb_dout0[31]
  PIN bb_dout0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 828.960 4.000 829.560 ;
    END
  END bb_dout0[3]
  PIN bb_dout0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 860.920 4.000 861.520 ;
    END
  END bb_dout0[4]
  PIN bb_dout0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 888.120 4.000 888.720 ;
    END
  END bb_dout0[5]
  PIN bb_dout0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 915.320 4.000 915.920 ;
    END
  END bb_dout0[6]
  PIN bb_dout0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 942.520 4.000 943.120 ;
    END
  END bb_dout0[7]
  PIN bb_dout0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 969.040 4.000 969.640 ;
    END
  END bb_dout0[8]
  PIN bb_dout0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 996.240 4.000 996.840 ;
    END
  END bb_dout0[9]
  PIN bb_dout1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 737.160 4.000 737.760 ;
    END
  END bb_dout1[0]
  PIN bb_dout1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1028.880 4.000 1029.480 ;
    END
  END bb_dout1[10]
  PIN bb_dout1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1056.080 4.000 1056.680 ;
    END
  END bb_dout1[11]
  PIN bb_dout1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1082.600 4.000 1083.200 ;
    END
  END bb_dout1[12]
  PIN bb_dout1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1109.800 4.000 1110.400 ;
    END
  END bb_dout1[13]
  PIN bb_dout1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1137.000 4.000 1137.600 ;
    END
  END bb_dout1[14]
  PIN bb_dout1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1164.200 4.000 1164.800 ;
    END
  END bb_dout1[15]
  PIN bb_dout1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1190.720 4.000 1191.320 ;
    END
  END bb_dout1[16]
  PIN bb_dout1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1217.920 4.000 1218.520 ;
    END
  END bb_dout1[17]
  PIN bb_dout1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1245.120 4.000 1245.720 ;
    END
  END bb_dout1[18]
  PIN bb_dout1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1272.320 4.000 1272.920 ;
    END
  END bb_dout1[19]
  PIN bb_dout1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 769.120 4.000 769.720 ;
    END
  END bb_dout1[1]
  PIN bb_dout1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1298.840 4.000 1299.440 ;
    END
  END bb_dout1[20]
  PIN bb_dout1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1326.040 4.000 1326.640 ;
    END
  END bb_dout1[21]
  PIN bb_dout1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1353.240 4.000 1353.840 ;
    END
  END bb_dout1[22]
  PIN bb_dout1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1380.440 4.000 1381.040 ;
    END
  END bb_dout1[23]
  PIN bb_dout1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1406.960 4.000 1407.560 ;
    END
  END bb_dout1[24]
  PIN bb_dout1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1434.160 4.000 1434.760 ;
    END
  END bb_dout1[25]
  PIN bb_dout1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1461.360 4.000 1461.960 ;
    END
  END bb_dout1[26]
  PIN bb_dout1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1488.560 4.000 1489.160 ;
    END
  END bb_dout1[27]
  PIN bb_dout1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1515.080 4.000 1515.680 ;
    END
  END bb_dout1[28]
  PIN bb_dout1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1542.280 4.000 1542.880 ;
    END
  END bb_dout1[29]
  PIN bb_dout1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 801.760 4.000 802.360 ;
    END
  END bb_dout1[2]
  PIN bb_dout1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1569.480 4.000 1570.080 ;
    END
  END bb_dout1[30]
  PIN bb_dout1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1596.680 4.000 1597.280 ;
    END
  END bb_dout1[31]
  PIN bb_dout1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 834.400 4.000 835.000 ;
    END
  END bb_dout1[3]
  PIN bb_dout1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 866.360 4.000 866.960 ;
    END
  END bb_dout1[4]
  PIN bb_dout1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 893.560 4.000 894.160 ;
    END
  END bb_dout1[5]
  PIN bb_dout1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 920.760 4.000 921.360 ;
    END
  END bb_dout1[6]
  PIN bb_dout1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 947.960 4.000 948.560 ;
    END
  END bb_dout1[7]
  PIN bb_dout1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 974.480 4.000 975.080 ;
    END
  END bb_dout1[8]
  PIN bb_dout1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1001.680 4.000 1002.280 ;
    END
  END bb_dout1[9]
  PIN bb_web0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 709.960 4.000 710.560 ;
    END
  END bb_web0
  PIN bb_wmask0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 742.600 4.000 743.200 ;
    END
  END bb_wmask0[0]
  PIN bb_wmask0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 774.560 4.000 775.160 ;
    END
  END bb_wmask0[1]
  PIN bb_wmask0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 807.200 4.000 807.800 ;
    END
  END bb_wmask0[2]
  PIN bb_wmask0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 839.840 4.000 840.440 ;
    END
  END bb_wmask0[3]
  PIN clk_g
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.670 0.000 10.950 4.000 ;
    END
  END clk_g
  PIN io_gecerli
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.770 0.000 96.050 4.000 ;
    END
  END io_gecerli
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.930 0.000 117.210 4.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 543.810 0.000 544.090 4.000 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 586.590 0.000 586.870 4.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 628.910 0.000 629.190 4.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 671.690 0.000 671.970 4.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 714.470 0.000 714.750 4.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 757.250 0.000 757.530 4.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 799.570 0.000 799.850 4.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 842.350 0.000 842.630 4.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 885.130 0.000 885.410 4.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 927.910 0.000 928.190 4.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.710 0.000 159.990 4.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 970.230 0.000 970.510 4.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1013.010 0.000 1013.290 4.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1055.790 0.000 1056.070 4.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1098.570 0.000 1098.850 4.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1140.890 0.000 1141.170 4.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1183.670 0.000 1183.950 4.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1226.450 0.000 1226.730 4.000 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1269.230 0.000 1269.510 4.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1311.550 0.000 1311.830 4.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1354.330 0.000 1354.610 4.000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.490 0.000 202.770 4.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1397.110 0.000 1397.390 4.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1439.890 0.000 1440.170 4.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1482.210 0.000 1482.490 4.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1503.830 0.000 1504.110 4.000 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1524.990 0.000 1525.270 4.000 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1546.150 0.000 1546.430 4.000 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1567.770 0.000 1568.050 4.000 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1588.930 0.000 1589.210 4.000 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 245.270 0.000 245.550 4.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.590 0.000 287.870 4.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 330.370 0.000 330.650 4.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 373.150 0.000 373.430 4.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.930 0.000 416.210 4.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 458.250 0.000 458.530 4.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 501.030 0.000 501.310 4.000 ;
    END
  END io_oeb[9]
  PIN io_ps[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.550 0.000 138.830 4.000 ;
    END
  END io_ps[0]
  PIN io_ps[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.970 0.000 565.250 4.000 ;
    END
  END io_ps[10]
  PIN io_ps[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 607.750 0.000 608.030 4.000 ;
    END
  END io_ps[11]
  PIN io_ps[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 650.530 0.000 650.810 4.000 ;
    END
  END io_ps[12]
  PIN io_ps[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 692.850 0.000 693.130 4.000 ;
    END
  END io_ps[13]
  PIN io_ps[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 735.630 0.000 735.910 4.000 ;
    END
  END io_ps[14]
  PIN io_ps[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 778.410 0.000 778.690 4.000 ;
    END
  END io_ps[15]
  PIN io_ps[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 821.190 0.000 821.470 4.000 ;
    END
  END io_ps[16]
  PIN io_ps[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 863.510 0.000 863.790 4.000 ;
    END
  END io_ps[17]
  PIN io_ps[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 906.290 0.000 906.570 4.000 ;
    END
  END io_ps[18]
  PIN io_ps[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 949.070 0.000 949.350 4.000 ;
    END
  END io_ps[19]
  PIN io_ps[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.870 0.000 181.150 4.000 ;
    END
  END io_ps[1]
  PIN io_ps[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 991.850 0.000 992.130 4.000 ;
    END
  END io_ps[20]
  PIN io_ps[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1034.170 0.000 1034.450 4.000 ;
    END
  END io_ps[21]
  PIN io_ps[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1076.950 0.000 1077.230 4.000 ;
    END
  END io_ps[22]
  PIN io_ps[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1119.730 0.000 1120.010 4.000 ;
    END
  END io_ps[23]
  PIN io_ps[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1162.510 0.000 1162.790 4.000 ;
    END
  END io_ps[24]
  PIN io_ps[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1204.830 0.000 1205.110 4.000 ;
    END
  END io_ps[25]
  PIN io_ps[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1247.610 0.000 1247.890 4.000 ;
    END
  END io_ps[26]
  PIN io_ps[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1290.390 0.000 1290.670 4.000 ;
    END
  END io_ps[27]
  PIN io_ps[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1333.170 0.000 1333.450 4.000 ;
    END
  END io_ps[28]
  PIN io_ps[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1375.490 0.000 1375.770 4.000 ;
    END
  END io_ps[29]
  PIN io_ps[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.650 0.000 223.930 4.000 ;
    END
  END io_ps[2]
  PIN io_ps[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1418.270 0.000 1418.550 4.000 ;
    END
  END io_ps[30]
  PIN io_ps[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1461.050 0.000 1461.330 4.000 ;
    END
  END io_ps[31]
  PIN io_ps[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.430 0.000 266.710 4.000 ;
    END
  END io_ps[3]
  PIN io_ps[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.210 0.000 309.490 4.000 ;
    END
  END io_ps[4]
  PIN io_ps[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.530 0.000 351.810 4.000 ;
    END
  END io_ps[5]
  PIN io_ps[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 394.310 0.000 394.590 4.000 ;
    END
  END io_ps[6]
  PIN io_ps[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 437.090 0.000 437.370 4.000 ;
    END
  END io_ps[7]
  PIN io_ps[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 479.870 0.000 480.150 4.000 ;
    END
  END io_ps[8]
  PIN io_ps[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 522.190 0.000 522.470 4.000 ;
    END
  END io_ps[9]
  PIN rst_g
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.830 0.000 32.110 4.000 ;
    END
  END rst_g
  PIN rx
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.610 0.000 74.890 4.000 ;
    END
  END rx
  PIN tx
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.990 0.000 53.270 4.000 ;
    END
  END tx
  PIN vb_addr0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.720 4.000 18.320 ;
    END
  END vb_addr0[0]
  PIN vb_addr0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 310.120 4.000 310.720 ;
    END
  END vb_addr0[10]
  PIN vb_addr0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 336.640 4.000 337.240 ;
    END
  END vb_addr0[11]
  PIN vb_addr0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 363.840 4.000 364.440 ;
    END
  END vb_addr0[12]
  PIN vb_addr0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 50.360 4.000 50.960 ;
    END
  END vb_addr0[1]
  PIN vb_addr0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.000 4.000 83.600 ;
    END
  END vb_addr0[2]
  PIN vb_addr0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 114.960 4.000 115.560 ;
    END
  END vb_addr0[3]
  PIN vb_addr0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 147.600 4.000 148.200 ;
    END
  END vb_addr0[4]
  PIN vb_addr0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 174.800 4.000 175.400 ;
    END
  END vb_addr0[5]
  PIN vb_addr0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 202.000 4.000 202.600 ;
    END
  END vb_addr0[6]
  PIN vb_addr0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 228.520 4.000 229.120 ;
    END
  END vb_addr0[7]
  PIN vb_addr0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 255.720 4.000 256.320 ;
    END
  END vb_addr0[8]
  PIN vb_addr0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 282.920 4.000 283.520 ;
    END
  END vb_addr0[9]
  PIN vb_addr1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.160 4.000 23.760 ;
    END
  END vb_addr1[0]
  PIN vb_addr1[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 315.560 4.000 316.160 ;
    END
  END vb_addr1[10]
  PIN vb_addr1[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 342.080 4.000 342.680 ;
    END
  END vb_addr1[11]
  PIN vb_addr1[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 369.280 4.000 369.880 ;
    END
  END vb_addr1[12]
  PIN vb_addr1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.800 4.000 56.400 ;
    END
  END vb_addr1[1]
  PIN vb_addr1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END vb_addr1[2]
  PIN vb_addr1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 120.400 4.000 121.000 ;
    END
  END vb_addr1[3]
  PIN vb_addr1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.040 4.000 153.640 ;
    END
  END vb_addr1[4]
  PIN vb_addr1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.240 4.000 180.840 ;
    END
  END vb_addr1[5]
  PIN vb_addr1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 207.440 4.000 208.040 ;
    END
  END vb_addr1[6]
  PIN vb_addr1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 233.960 4.000 234.560 ;
    END
  END vb_addr1[7]
  PIN vb_addr1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 261.160 4.000 261.760 ;
    END
  END vb_addr1[8]
  PIN vb_addr1[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 288.360 4.000 288.960 ;
    END
  END vb_addr1[9]
  PIN vb_csb0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.080 4.000 2.680 ;
    END
  END vb_csb0
  PIN vb_csb1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END vb_csb1
  PIN vb_din0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 28.600 4.000 29.200 ;
    END
  END vb_din0[0]
  PIN vb_din0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 321.000 4.000 321.600 ;
    END
  END vb_din0[10]
  PIN vb_din0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 347.520 4.000 348.120 ;
    END
  END vb_din0[11]
  PIN vb_din0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 374.720 4.000 375.320 ;
    END
  END vb_din0[12]
  PIN vb_din0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 391.040 4.000 391.640 ;
    END
  END vb_din0[13]
  PIN vb_din0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 407.360 4.000 407.960 ;
    END
  END vb_din0[14]
  PIN vb_din0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 423.680 4.000 424.280 ;
    END
  END vb_din0[15]
  PIN vb_din0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 439.320 4.000 439.920 ;
    END
  END vb_din0[16]
  PIN vb_din0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 455.640 4.000 456.240 ;
    END
  END vb_din0[17]
  PIN vb_din0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 471.960 4.000 472.560 ;
    END
  END vb_din0[18]
  PIN vb_din0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 488.280 4.000 488.880 ;
    END
  END vb_din0[19]
  PIN vb_din0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END vb_din0[1]
  PIN vb_din0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 504.600 4.000 505.200 ;
    END
  END vb_din0[20]
  PIN vb_din0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 520.920 4.000 521.520 ;
    END
  END vb_din0[21]
  PIN vb_din0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 536.560 4.000 537.160 ;
    END
  END vb_din0[22]
  PIN vb_din0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 552.880 4.000 553.480 ;
    END
  END vb_din0[23]
  PIN vb_din0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 569.200 4.000 569.800 ;
    END
  END vb_din0[24]
  PIN vb_din0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 585.520 4.000 586.120 ;
    END
  END vb_din0[25]
  PIN vb_din0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 601.840 4.000 602.440 ;
    END
  END vb_din0[26]
  PIN vb_din0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 618.160 4.000 618.760 ;
    END
  END vb_din0[27]
  PIN vb_din0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 634.480 4.000 635.080 ;
    END
  END vb_din0[28]
  PIN vb_din0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 650.120 4.000 650.720 ;
    END
  END vb_din0[29]
  PIN vb_din0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.880 4.000 94.480 ;
    END
  END vb_din0[2]
  PIN vb_din0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 666.440 4.000 667.040 ;
    END
  END vb_din0[30]
  PIN vb_din0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 682.760 4.000 683.360 ;
    END
  END vb_din0[31]
  PIN vb_din0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.840 4.000 126.440 ;
    END
  END vb_din0[3]
  PIN vb_din0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 158.480 4.000 159.080 ;
    END
  END vb_din0[4]
  PIN vb_din0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 185.680 4.000 186.280 ;
    END
  END vb_din0[5]
  PIN vb_din0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 212.880 4.000 213.480 ;
    END
  END vb_din0[6]
  PIN vb_din0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 239.400 4.000 240.000 ;
    END
  END vb_din0[7]
  PIN vb_din0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 266.600 4.000 267.200 ;
    END
  END vb_din0[8]
  PIN vb_din0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 293.800 4.000 294.400 ;
    END
  END vb_din0[9]
  PIN vb_dout0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END vb_dout0[0]
  PIN vb_dout0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 325.760 4.000 326.360 ;
    END
  END vb_dout0[10]
  PIN vb_dout0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 352.960 4.000 353.560 ;
    END
  END vb_dout0[11]
  PIN vb_dout0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 380.160 4.000 380.760 ;
    END
  END vb_dout0[12]
  PIN vb_dout0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 396.480 4.000 397.080 ;
    END
  END vb_dout0[13]
  PIN vb_dout0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 412.800 4.000 413.400 ;
    END
  END vb_dout0[14]
  PIN vb_dout0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 428.440 4.000 429.040 ;
    END
  END vb_dout0[15]
  PIN vb_dout0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 444.760 4.000 445.360 ;
    END
  END vb_dout0[16]
  PIN vb_dout0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 461.080 4.000 461.680 ;
    END
  END vb_dout0[17]
  PIN vb_dout0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 477.400 4.000 478.000 ;
    END
  END vb_dout0[18]
  PIN vb_dout0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 493.720 4.000 494.320 ;
    END
  END vb_dout0[19]
  PIN vb_dout0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.680 4.000 67.280 ;
    END
  END vb_dout0[1]
  PIN vb_dout0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 510.040 4.000 510.640 ;
    END
  END vb_dout0[20]
  PIN vb_dout0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 526.360 4.000 526.960 ;
    END
  END vb_dout0[21]
  PIN vb_dout0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 542.000 4.000 542.600 ;
    END
  END vb_dout0[22]
  PIN vb_dout0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 558.320 4.000 558.920 ;
    END
  END vb_dout0[23]
  PIN vb_dout0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 574.640 4.000 575.240 ;
    END
  END vb_dout0[24]
  PIN vb_dout0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 590.960 4.000 591.560 ;
    END
  END vb_dout0[25]
  PIN vb_dout0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 607.280 4.000 607.880 ;
    END
  END vb_dout0[26]
  PIN vb_dout0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 623.600 4.000 624.200 ;
    END
  END vb_dout0[27]
  PIN vb_dout0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 639.920 4.000 640.520 ;
    END
  END vb_dout0[28]
  PIN vb_dout0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 655.560 4.000 656.160 ;
    END
  END vb_dout0[29]
  PIN vb_dout0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 99.320 4.000 99.920 ;
    END
  END vb_dout0[2]
  PIN vb_dout0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 671.880 4.000 672.480 ;
    END
  END vb_dout0[30]
  PIN vb_dout0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 688.200 4.000 688.800 ;
    END
  END vb_dout0[31]
  PIN vb_dout0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 131.280 4.000 131.880 ;
    END
  END vb_dout0[3]
  PIN vb_dout0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.920 4.000 164.520 ;
    END
  END vb_dout0[4]
  PIN vb_dout0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 191.120 4.000 191.720 ;
    END
  END vb_dout0[5]
  PIN vb_dout0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 217.640 4.000 218.240 ;
    END
  END vb_dout0[6]
  PIN vb_dout0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 244.840 4.000 245.440 ;
    END
  END vb_dout0[7]
  PIN vb_dout0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 272.040 4.000 272.640 ;
    END
  END vb_dout0[8]
  PIN vb_dout0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 299.240 4.000 299.840 ;
    END
  END vb_dout0[9]
  PIN vb_dout1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 39.480 4.000 40.080 ;
    END
  END vb_dout1[0]
  PIN vb_dout1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 331.200 4.000 331.800 ;
    END
  END vb_dout1[10]
  PIN vb_dout1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 358.400 4.000 359.000 ;
    END
  END vb_dout1[11]
  PIN vb_dout1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 385.600 4.000 386.200 ;
    END
  END vb_dout1[12]
  PIN vb_dout1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 401.920 4.000 402.520 ;
    END
  END vb_dout1[13]
  PIN vb_dout1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 418.240 4.000 418.840 ;
    END
  END vb_dout1[14]
  PIN vb_dout1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 433.880 4.000 434.480 ;
    END
  END vb_dout1[15]
  PIN vb_dout1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 450.200 4.000 450.800 ;
    END
  END vb_dout1[16]
  PIN vb_dout1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 466.520 4.000 467.120 ;
    END
  END vb_dout1[17]
  PIN vb_dout1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 482.840 4.000 483.440 ;
    END
  END vb_dout1[18]
  PIN vb_dout1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 499.160 4.000 499.760 ;
    END
  END vb_dout1[19]
  PIN vb_dout1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.120 4.000 72.720 ;
    END
  END vb_dout1[1]
  PIN vb_dout1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 515.480 4.000 516.080 ;
    END
  END vb_dout1[20]
  PIN vb_dout1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 531.800 4.000 532.400 ;
    END
  END vb_dout1[21]
  PIN vb_dout1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 547.440 4.000 548.040 ;
    END
  END vb_dout1[22]
  PIN vb_dout1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 563.760 4.000 564.360 ;
    END
  END vb_dout1[23]
  PIN vb_dout1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 580.080 4.000 580.680 ;
    END
  END vb_dout1[24]
  PIN vb_dout1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 596.400 4.000 597.000 ;
    END
  END vb_dout1[25]
  PIN vb_dout1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 612.720 4.000 613.320 ;
    END
  END vb_dout1[26]
  PIN vb_dout1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 629.040 4.000 629.640 ;
    END
  END vb_dout1[27]
  PIN vb_dout1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 644.680 4.000 645.280 ;
    END
  END vb_dout1[28]
  PIN vb_dout1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 661.000 4.000 661.600 ;
    END
  END vb_dout1[29]
  PIN vb_dout1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 104.760 4.000 105.360 ;
    END
  END vb_dout1[2]
  PIN vb_dout1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 677.320 4.000 677.920 ;
    END
  END vb_dout1[30]
  PIN vb_dout1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 693.640 4.000 694.240 ;
    END
  END vb_dout1[31]
  PIN vb_dout1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.720 4.000 137.320 ;
    END
  END vb_dout1[3]
  PIN vb_dout1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 169.360 4.000 169.960 ;
    END
  END vb_dout1[4]
  PIN vb_dout1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 196.560 4.000 197.160 ;
    END
  END vb_dout1[5]
  PIN vb_dout1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 223.080 4.000 223.680 ;
    END
  END vb_dout1[6]
  PIN vb_dout1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 250.280 4.000 250.880 ;
    END
  END vb_dout1[7]
  PIN vb_dout1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 277.480 4.000 278.080 ;
    END
  END vb_dout1[8]
  PIN vb_dout1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 304.680 4.000 305.280 ;
    END
  END vb_dout1[9]
  PIN vb_web0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.280 4.000 12.880 ;
    END
  END vb_web0
  PIN vb_wmask0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.920 4.000 45.520 ;
    END
  END vb_wmask0[0]
  PIN vb_wmask0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 77.560 4.000 78.160 ;
    END
  END vb_wmask0[1]
  PIN vb_wmask0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 109.520 4.000 110.120 ;
    END
  END vb_wmask0[2]
  PIN vb_wmask0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.160 4.000 142.760 ;
    END
  END vb_wmask0[3]
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.840 10.640 1251.440 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1403.440 10.640 1405.040 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1557.040 10.640 1558.640 1588.720 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1326.640 10.640 1328.240 1588.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 1480.240 10.640 1481.840 1588.720 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 1594.360 1588.565 ;
      LAYER met1 ;
        RECT 1.910 9.900 1594.360 1588.720 ;
      LAYER met2 ;
        RECT 1.940 4.280 1589.200 1597.165 ;
        RECT 1.940 2.195 10.390 4.280 ;
        RECT 11.230 2.195 31.550 4.280 ;
        RECT 32.390 2.195 52.710 4.280 ;
        RECT 53.550 2.195 74.330 4.280 ;
        RECT 75.170 2.195 95.490 4.280 ;
        RECT 96.330 2.195 116.650 4.280 ;
        RECT 117.490 2.195 138.270 4.280 ;
        RECT 139.110 2.195 159.430 4.280 ;
        RECT 160.270 2.195 180.590 4.280 ;
        RECT 181.430 2.195 202.210 4.280 ;
        RECT 203.050 2.195 223.370 4.280 ;
        RECT 224.210 2.195 244.990 4.280 ;
        RECT 245.830 2.195 266.150 4.280 ;
        RECT 266.990 2.195 287.310 4.280 ;
        RECT 288.150 2.195 308.930 4.280 ;
        RECT 309.770 2.195 330.090 4.280 ;
        RECT 330.930 2.195 351.250 4.280 ;
        RECT 352.090 2.195 372.870 4.280 ;
        RECT 373.710 2.195 394.030 4.280 ;
        RECT 394.870 2.195 415.650 4.280 ;
        RECT 416.490 2.195 436.810 4.280 ;
        RECT 437.650 2.195 457.970 4.280 ;
        RECT 458.810 2.195 479.590 4.280 ;
        RECT 480.430 2.195 500.750 4.280 ;
        RECT 501.590 2.195 521.910 4.280 ;
        RECT 522.750 2.195 543.530 4.280 ;
        RECT 544.370 2.195 564.690 4.280 ;
        RECT 565.530 2.195 586.310 4.280 ;
        RECT 587.150 2.195 607.470 4.280 ;
        RECT 608.310 2.195 628.630 4.280 ;
        RECT 629.470 2.195 650.250 4.280 ;
        RECT 651.090 2.195 671.410 4.280 ;
        RECT 672.250 2.195 692.570 4.280 ;
        RECT 693.410 2.195 714.190 4.280 ;
        RECT 715.030 2.195 735.350 4.280 ;
        RECT 736.190 2.195 756.970 4.280 ;
        RECT 757.810 2.195 778.130 4.280 ;
        RECT 778.970 2.195 799.290 4.280 ;
        RECT 800.130 2.195 820.910 4.280 ;
        RECT 821.750 2.195 842.070 4.280 ;
        RECT 842.910 2.195 863.230 4.280 ;
        RECT 864.070 2.195 884.850 4.280 ;
        RECT 885.690 2.195 906.010 4.280 ;
        RECT 906.850 2.195 927.630 4.280 ;
        RECT 928.470 2.195 948.790 4.280 ;
        RECT 949.630 2.195 969.950 4.280 ;
        RECT 970.790 2.195 991.570 4.280 ;
        RECT 992.410 2.195 1012.730 4.280 ;
        RECT 1013.570 2.195 1033.890 4.280 ;
        RECT 1034.730 2.195 1055.510 4.280 ;
        RECT 1056.350 2.195 1076.670 4.280 ;
        RECT 1077.510 2.195 1098.290 4.280 ;
        RECT 1099.130 2.195 1119.450 4.280 ;
        RECT 1120.290 2.195 1140.610 4.280 ;
        RECT 1141.450 2.195 1162.230 4.280 ;
        RECT 1163.070 2.195 1183.390 4.280 ;
        RECT 1184.230 2.195 1204.550 4.280 ;
        RECT 1205.390 2.195 1226.170 4.280 ;
        RECT 1227.010 2.195 1247.330 4.280 ;
        RECT 1248.170 2.195 1268.950 4.280 ;
        RECT 1269.790 2.195 1290.110 4.280 ;
        RECT 1290.950 2.195 1311.270 4.280 ;
        RECT 1312.110 2.195 1332.890 4.280 ;
        RECT 1333.730 2.195 1354.050 4.280 ;
        RECT 1354.890 2.195 1375.210 4.280 ;
        RECT 1376.050 2.195 1396.830 4.280 ;
        RECT 1397.670 2.195 1417.990 4.280 ;
        RECT 1418.830 2.195 1439.610 4.280 ;
        RECT 1440.450 2.195 1460.770 4.280 ;
        RECT 1461.610 2.195 1481.930 4.280 ;
        RECT 1482.770 2.195 1503.550 4.280 ;
        RECT 1504.390 2.195 1524.710 4.280 ;
        RECT 1525.550 2.195 1545.870 4.280 ;
        RECT 1546.710 2.195 1567.490 4.280 ;
        RECT 1568.330 2.195 1588.650 4.280 ;
      LAYER met3 ;
        RECT 4.400 1596.280 1558.640 1597.145 ;
        RECT 4.000 1592.240 1558.640 1596.280 ;
        RECT 4.400 1590.840 1558.640 1592.240 ;
        RECT 4.000 1586.800 1558.640 1590.840 ;
        RECT 4.400 1585.400 1558.640 1586.800 ;
        RECT 4.000 1581.360 1558.640 1585.400 ;
        RECT 4.400 1579.960 1558.640 1581.360 ;
        RECT 4.000 1575.920 1558.640 1579.960 ;
        RECT 4.400 1574.520 1558.640 1575.920 ;
        RECT 4.000 1570.480 1558.640 1574.520 ;
        RECT 4.400 1569.080 1558.640 1570.480 ;
        RECT 4.000 1565.040 1558.640 1569.080 ;
        RECT 4.400 1563.640 1558.640 1565.040 ;
        RECT 4.000 1559.600 1558.640 1563.640 ;
        RECT 4.400 1558.200 1558.640 1559.600 ;
        RECT 4.000 1554.160 1558.640 1558.200 ;
        RECT 4.400 1552.760 1558.640 1554.160 ;
        RECT 4.000 1548.720 1558.640 1552.760 ;
        RECT 4.400 1547.320 1558.640 1548.720 ;
        RECT 4.000 1543.280 1558.640 1547.320 ;
        RECT 4.400 1541.880 1558.640 1543.280 ;
        RECT 4.000 1537.840 1558.640 1541.880 ;
        RECT 4.400 1536.440 1558.640 1537.840 ;
        RECT 4.000 1532.400 1558.640 1536.440 ;
        RECT 4.400 1531.000 1558.640 1532.400 ;
        RECT 4.000 1526.960 1558.640 1531.000 ;
        RECT 4.400 1525.560 1558.640 1526.960 ;
        RECT 4.000 1521.520 1558.640 1525.560 ;
        RECT 4.400 1520.120 1558.640 1521.520 ;
        RECT 4.000 1516.080 1558.640 1520.120 ;
        RECT 4.400 1514.680 1558.640 1516.080 ;
        RECT 4.000 1510.640 1558.640 1514.680 ;
        RECT 4.400 1509.240 1558.640 1510.640 ;
        RECT 4.000 1505.200 1558.640 1509.240 ;
        RECT 4.400 1503.800 1558.640 1505.200 ;
        RECT 4.000 1499.760 1558.640 1503.800 ;
        RECT 4.400 1498.360 1558.640 1499.760 ;
        RECT 4.000 1495.000 1558.640 1498.360 ;
        RECT 4.400 1493.600 1558.640 1495.000 ;
        RECT 4.000 1489.560 1558.640 1493.600 ;
        RECT 4.400 1488.160 1558.640 1489.560 ;
        RECT 4.000 1484.120 1558.640 1488.160 ;
        RECT 4.400 1482.720 1558.640 1484.120 ;
        RECT 4.000 1478.680 1558.640 1482.720 ;
        RECT 4.400 1477.280 1558.640 1478.680 ;
        RECT 4.000 1473.240 1558.640 1477.280 ;
        RECT 4.400 1471.840 1558.640 1473.240 ;
        RECT 4.000 1467.800 1558.640 1471.840 ;
        RECT 4.400 1466.400 1558.640 1467.800 ;
        RECT 4.000 1462.360 1558.640 1466.400 ;
        RECT 4.400 1460.960 1558.640 1462.360 ;
        RECT 4.000 1456.920 1558.640 1460.960 ;
        RECT 4.400 1455.520 1558.640 1456.920 ;
        RECT 4.000 1451.480 1558.640 1455.520 ;
        RECT 4.400 1450.080 1558.640 1451.480 ;
        RECT 4.000 1446.040 1558.640 1450.080 ;
        RECT 4.400 1444.640 1558.640 1446.040 ;
        RECT 4.000 1440.600 1558.640 1444.640 ;
        RECT 4.400 1439.200 1558.640 1440.600 ;
        RECT 4.000 1435.160 1558.640 1439.200 ;
        RECT 4.400 1433.760 1558.640 1435.160 ;
        RECT 4.000 1429.720 1558.640 1433.760 ;
        RECT 4.400 1428.320 1558.640 1429.720 ;
        RECT 4.000 1424.280 1558.640 1428.320 ;
        RECT 4.400 1422.880 1558.640 1424.280 ;
        RECT 4.000 1418.840 1558.640 1422.880 ;
        RECT 4.400 1417.440 1558.640 1418.840 ;
        RECT 4.000 1413.400 1558.640 1417.440 ;
        RECT 4.400 1412.000 1558.640 1413.400 ;
        RECT 4.000 1407.960 1558.640 1412.000 ;
        RECT 4.400 1406.560 1558.640 1407.960 ;
        RECT 4.000 1402.520 1558.640 1406.560 ;
        RECT 4.400 1401.120 1558.640 1402.520 ;
        RECT 4.000 1397.080 1558.640 1401.120 ;
        RECT 4.400 1395.680 1558.640 1397.080 ;
        RECT 4.000 1391.640 1558.640 1395.680 ;
        RECT 4.400 1390.240 1558.640 1391.640 ;
        RECT 4.000 1386.880 1558.640 1390.240 ;
        RECT 4.400 1385.480 1558.640 1386.880 ;
        RECT 4.000 1381.440 1558.640 1385.480 ;
        RECT 4.400 1380.040 1558.640 1381.440 ;
        RECT 4.000 1376.000 1558.640 1380.040 ;
        RECT 4.400 1374.600 1558.640 1376.000 ;
        RECT 4.000 1370.560 1558.640 1374.600 ;
        RECT 4.400 1369.160 1558.640 1370.560 ;
        RECT 4.000 1365.120 1558.640 1369.160 ;
        RECT 4.400 1363.720 1558.640 1365.120 ;
        RECT 4.000 1359.680 1558.640 1363.720 ;
        RECT 4.400 1358.280 1558.640 1359.680 ;
        RECT 4.000 1354.240 1558.640 1358.280 ;
        RECT 4.400 1352.840 1558.640 1354.240 ;
        RECT 4.000 1348.800 1558.640 1352.840 ;
        RECT 4.400 1347.400 1558.640 1348.800 ;
        RECT 4.000 1343.360 1558.640 1347.400 ;
        RECT 4.400 1341.960 1558.640 1343.360 ;
        RECT 4.000 1337.920 1558.640 1341.960 ;
        RECT 4.400 1336.520 1558.640 1337.920 ;
        RECT 4.000 1332.480 1558.640 1336.520 ;
        RECT 4.400 1331.080 1558.640 1332.480 ;
        RECT 4.000 1327.040 1558.640 1331.080 ;
        RECT 4.400 1325.640 1558.640 1327.040 ;
        RECT 4.000 1321.600 1558.640 1325.640 ;
        RECT 4.400 1320.200 1558.640 1321.600 ;
        RECT 4.000 1316.160 1558.640 1320.200 ;
        RECT 4.400 1314.760 1558.640 1316.160 ;
        RECT 4.000 1310.720 1558.640 1314.760 ;
        RECT 4.400 1309.320 1558.640 1310.720 ;
        RECT 4.000 1305.280 1558.640 1309.320 ;
        RECT 4.400 1303.880 1558.640 1305.280 ;
        RECT 4.000 1299.840 1558.640 1303.880 ;
        RECT 4.400 1298.440 1558.640 1299.840 ;
        RECT 4.000 1294.400 1558.640 1298.440 ;
        RECT 4.400 1293.000 1558.640 1294.400 ;
        RECT 4.000 1288.960 1558.640 1293.000 ;
        RECT 4.400 1287.560 1558.640 1288.960 ;
        RECT 4.000 1283.520 1558.640 1287.560 ;
        RECT 4.400 1282.120 1558.640 1283.520 ;
        RECT 4.000 1278.760 1558.640 1282.120 ;
        RECT 4.400 1277.360 1558.640 1278.760 ;
        RECT 4.000 1273.320 1558.640 1277.360 ;
        RECT 4.400 1271.920 1558.640 1273.320 ;
        RECT 4.000 1267.880 1558.640 1271.920 ;
        RECT 4.400 1266.480 1558.640 1267.880 ;
        RECT 4.000 1262.440 1558.640 1266.480 ;
        RECT 4.400 1261.040 1558.640 1262.440 ;
        RECT 4.000 1257.000 1558.640 1261.040 ;
        RECT 4.400 1255.600 1558.640 1257.000 ;
        RECT 4.000 1251.560 1558.640 1255.600 ;
        RECT 4.400 1250.160 1558.640 1251.560 ;
        RECT 4.000 1246.120 1558.640 1250.160 ;
        RECT 4.400 1244.720 1558.640 1246.120 ;
        RECT 4.000 1240.680 1558.640 1244.720 ;
        RECT 4.400 1239.280 1558.640 1240.680 ;
        RECT 4.000 1235.240 1558.640 1239.280 ;
        RECT 4.400 1233.840 1558.640 1235.240 ;
        RECT 4.000 1229.800 1558.640 1233.840 ;
        RECT 4.400 1228.400 1558.640 1229.800 ;
        RECT 4.000 1224.360 1558.640 1228.400 ;
        RECT 4.400 1222.960 1558.640 1224.360 ;
        RECT 4.000 1218.920 1558.640 1222.960 ;
        RECT 4.400 1217.520 1558.640 1218.920 ;
        RECT 4.000 1213.480 1558.640 1217.520 ;
        RECT 4.400 1212.080 1558.640 1213.480 ;
        RECT 4.000 1208.040 1558.640 1212.080 ;
        RECT 4.400 1206.640 1558.640 1208.040 ;
        RECT 4.000 1202.600 1558.640 1206.640 ;
        RECT 4.400 1201.200 1558.640 1202.600 ;
        RECT 4.000 1197.160 1558.640 1201.200 ;
        RECT 4.400 1195.760 1558.640 1197.160 ;
        RECT 4.000 1191.720 1558.640 1195.760 ;
        RECT 4.400 1190.320 1558.640 1191.720 ;
        RECT 4.000 1186.280 1558.640 1190.320 ;
        RECT 4.400 1184.880 1558.640 1186.280 ;
        RECT 4.000 1180.840 1558.640 1184.880 ;
        RECT 4.400 1179.440 1558.640 1180.840 ;
        RECT 4.000 1176.080 1558.640 1179.440 ;
        RECT 4.400 1174.680 1558.640 1176.080 ;
        RECT 4.000 1170.640 1558.640 1174.680 ;
        RECT 4.400 1169.240 1558.640 1170.640 ;
        RECT 4.000 1165.200 1558.640 1169.240 ;
        RECT 4.400 1163.800 1558.640 1165.200 ;
        RECT 4.000 1159.760 1558.640 1163.800 ;
        RECT 4.400 1158.360 1558.640 1159.760 ;
        RECT 4.000 1154.320 1558.640 1158.360 ;
        RECT 4.400 1152.920 1558.640 1154.320 ;
        RECT 4.000 1148.880 1558.640 1152.920 ;
        RECT 4.400 1147.480 1558.640 1148.880 ;
        RECT 4.000 1143.440 1558.640 1147.480 ;
        RECT 4.400 1142.040 1558.640 1143.440 ;
        RECT 4.000 1138.000 1558.640 1142.040 ;
        RECT 4.400 1136.600 1558.640 1138.000 ;
        RECT 4.000 1132.560 1558.640 1136.600 ;
        RECT 4.400 1131.160 1558.640 1132.560 ;
        RECT 4.000 1127.120 1558.640 1131.160 ;
        RECT 4.400 1125.720 1558.640 1127.120 ;
        RECT 4.000 1121.680 1558.640 1125.720 ;
        RECT 4.400 1120.280 1558.640 1121.680 ;
        RECT 4.000 1116.240 1558.640 1120.280 ;
        RECT 4.400 1114.840 1558.640 1116.240 ;
        RECT 4.000 1110.800 1558.640 1114.840 ;
        RECT 4.400 1109.400 1558.640 1110.800 ;
        RECT 4.000 1105.360 1558.640 1109.400 ;
        RECT 4.400 1103.960 1558.640 1105.360 ;
        RECT 4.000 1099.920 1558.640 1103.960 ;
        RECT 4.400 1098.520 1558.640 1099.920 ;
        RECT 4.000 1094.480 1558.640 1098.520 ;
        RECT 4.400 1093.080 1558.640 1094.480 ;
        RECT 4.000 1089.040 1558.640 1093.080 ;
        RECT 4.400 1087.640 1558.640 1089.040 ;
        RECT 4.000 1083.600 1558.640 1087.640 ;
        RECT 4.400 1082.200 1558.640 1083.600 ;
        RECT 4.000 1078.160 1558.640 1082.200 ;
        RECT 4.400 1076.760 1558.640 1078.160 ;
        RECT 4.000 1072.720 1558.640 1076.760 ;
        RECT 4.400 1071.320 1558.640 1072.720 ;
        RECT 4.000 1067.960 1558.640 1071.320 ;
        RECT 4.400 1066.560 1558.640 1067.960 ;
        RECT 4.000 1062.520 1558.640 1066.560 ;
        RECT 4.400 1061.120 1558.640 1062.520 ;
        RECT 4.000 1057.080 1558.640 1061.120 ;
        RECT 4.400 1055.680 1558.640 1057.080 ;
        RECT 4.000 1051.640 1558.640 1055.680 ;
        RECT 4.400 1050.240 1558.640 1051.640 ;
        RECT 4.000 1046.200 1558.640 1050.240 ;
        RECT 4.400 1044.800 1558.640 1046.200 ;
        RECT 4.000 1040.760 1558.640 1044.800 ;
        RECT 4.400 1039.360 1558.640 1040.760 ;
        RECT 4.000 1035.320 1558.640 1039.360 ;
        RECT 4.400 1033.920 1558.640 1035.320 ;
        RECT 4.000 1029.880 1558.640 1033.920 ;
        RECT 4.400 1028.480 1558.640 1029.880 ;
        RECT 4.000 1024.440 1558.640 1028.480 ;
        RECT 4.400 1023.040 1558.640 1024.440 ;
        RECT 4.000 1019.000 1558.640 1023.040 ;
        RECT 4.400 1017.600 1558.640 1019.000 ;
        RECT 4.000 1013.560 1558.640 1017.600 ;
        RECT 4.400 1012.160 1558.640 1013.560 ;
        RECT 4.000 1008.120 1558.640 1012.160 ;
        RECT 4.400 1006.720 1558.640 1008.120 ;
        RECT 4.000 1002.680 1558.640 1006.720 ;
        RECT 4.400 1001.280 1558.640 1002.680 ;
        RECT 4.000 997.240 1558.640 1001.280 ;
        RECT 4.400 995.840 1558.640 997.240 ;
        RECT 4.000 991.800 1558.640 995.840 ;
        RECT 4.400 990.400 1558.640 991.800 ;
        RECT 4.000 986.360 1558.640 990.400 ;
        RECT 4.400 984.960 1558.640 986.360 ;
        RECT 4.000 980.920 1558.640 984.960 ;
        RECT 4.400 979.520 1558.640 980.920 ;
        RECT 4.000 975.480 1558.640 979.520 ;
        RECT 4.400 974.080 1558.640 975.480 ;
        RECT 4.000 970.040 1558.640 974.080 ;
        RECT 4.400 968.640 1558.640 970.040 ;
        RECT 4.000 964.600 1558.640 968.640 ;
        RECT 4.400 963.200 1558.640 964.600 ;
        RECT 4.000 959.840 1558.640 963.200 ;
        RECT 4.400 958.440 1558.640 959.840 ;
        RECT 4.000 954.400 1558.640 958.440 ;
        RECT 4.400 953.000 1558.640 954.400 ;
        RECT 4.000 948.960 1558.640 953.000 ;
        RECT 4.400 947.560 1558.640 948.960 ;
        RECT 4.000 943.520 1558.640 947.560 ;
        RECT 4.400 942.120 1558.640 943.520 ;
        RECT 4.000 938.080 1558.640 942.120 ;
        RECT 4.400 936.680 1558.640 938.080 ;
        RECT 4.000 932.640 1558.640 936.680 ;
        RECT 4.400 931.240 1558.640 932.640 ;
        RECT 4.000 927.200 1558.640 931.240 ;
        RECT 4.400 925.800 1558.640 927.200 ;
        RECT 4.000 921.760 1558.640 925.800 ;
        RECT 4.400 920.360 1558.640 921.760 ;
        RECT 4.000 916.320 1558.640 920.360 ;
        RECT 4.400 914.920 1558.640 916.320 ;
        RECT 4.000 910.880 1558.640 914.920 ;
        RECT 4.400 909.480 1558.640 910.880 ;
        RECT 4.000 905.440 1558.640 909.480 ;
        RECT 4.400 904.040 1558.640 905.440 ;
        RECT 4.000 900.000 1558.640 904.040 ;
        RECT 4.400 898.600 1558.640 900.000 ;
        RECT 4.000 894.560 1558.640 898.600 ;
        RECT 4.400 893.160 1558.640 894.560 ;
        RECT 4.000 889.120 1558.640 893.160 ;
        RECT 4.400 887.720 1558.640 889.120 ;
        RECT 4.000 883.680 1558.640 887.720 ;
        RECT 4.400 882.280 1558.640 883.680 ;
        RECT 4.000 878.240 1558.640 882.280 ;
        RECT 4.400 876.840 1558.640 878.240 ;
        RECT 4.000 872.800 1558.640 876.840 ;
        RECT 4.400 871.400 1558.640 872.800 ;
        RECT 4.000 867.360 1558.640 871.400 ;
        RECT 4.400 865.960 1558.640 867.360 ;
        RECT 4.000 861.920 1558.640 865.960 ;
        RECT 4.400 860.520 1558.640 861.920 ;
        RECT 4.000 856.480 1558.640 860.520 ;
        RECT 4.400 855.080 1558.640 856.480 ;
        RECT 4.000 851.720 1558.640 855.080 ;
        RECT 4.400 850.320 1558.640 851.720 ;
        RECT 4.000 846.280 1558.640 850.320 ;
        RECT 4.400 844.880 1558.640 846.280 ;
        RECT 4.000 840.840 1558.640 844.880 ;
        RECT 4.400 839.440 1558.640 840.840 ;
        RECT 4.000 835.400 1558.640 839.440 ;
        RECT 4.400 834.000 1558.640 835.400 ;
        RECT 4.000 829.960 1558.640 834.000 ;
        RECT 4.400 828.560 1558.640 829.960 ;
        RECT 4.000 824.520 1558.640 828.560 ;
        RECT 4.400 823.120 1558.640 824.520 ;
        RECT 4.000 819.080 1558.640 823.120 ;
        RECT 4.400 817.680 1558.640 819.080 ;
        RECT 4.000 813.640 1558.640 817.680 ;
        RECT 4.400 812.240 1558.640 813.640 ;
        RECT 4.000 808.200 1558.640 812.240 ;
        RECT 4.400 806.800 1558.640 808.200 ;
        RECT 4.000 802.760 1558.640 806.800 ;
        RECT 4.400 801.360 1558.640 802.760 ;
        RECT 4.000 797.320 1558.640 801.360 ;
        RECT 4.400 795.920 1558.640 797.320 ;
        RECT 4.000 791.880 1558.640 795.920 ;
        RECT 4.400 790.480 1558.640 791.880 ;
        RECT 4.000 786.440 1558.640 790.480 ;
        RECT 4.400 785.040 1558.640 786.440 ;
        RECT 4.000 781.000 1558.640 785.040 ;
        RECT 4.400 779.600 1558.640 781.000 ;
        RECT 4.000 775.560 1558.640 779.600 ;
        RECT 4.400 774.160 1558.640 775.560 ;
        RECT 4.000 770.120 1558.640 774.160 ;
        RECT 4.400 768.720 1558.640 770.120 ;
        RECT 4.000 764.680 1558.640 768.720 ;
        RECT 4.400 763.280 1558.640 764.680 ;
        RECT 4.000 759.240 1558.640 763.280 ;
        RECT 4.400 757.840 1558.640 759.240 ;
        RECT 4.000 753.800 1558.640 757.840 ;
        RECT 4.400 752.400 1558.640 753.800 ;
        RECT 4.000 749.040 1558.640 752.400 ;
        RECT 4.400 747.640 1558.640 749.040 ;
        RECT 4.000 743.600 1558.640 747.640 ;
        RECT 4.400 742.200 1558.640 743.600 ;
        RECT 4.000 738.160 1558.640 742.200 ;
        RECT 4.400 736.760 1558.640 738.160 ;
        RECT 4.000 732.720 1558.640 736.760 ;
        RECT 4.400 731.320 1558.640 732.720 ;
        RECT 4.000 727.280 1558.640 731.320 ;
        RECT 4.400 725.880 1558.640 727.280 ;
        RECT 4.000 721.840 1558.640 725.880 ;
        RECT 4.400 720.440 1558.640 721.840 ;
        RECT 4.000 716.400 1558.640 720.440 ;
        RECT 4.400 715.000 1558.640 716.400 ;
        RECT 4.000 710.960 1558.640 715.000 ;
        RECT 4.400 709.560 1558.640 710.960 ;
        RECT 4.000 705.520 1558.640 709.560 ;
        RECT 4.400 704.120 1558.640 705.520 ;
        RECT 4.000 700.080 1558.640 704.120 ;
        RECT 4.400 698.680 1558.640 700.080 ;
        RECT 4.000 694.640 1558.640 698.680 ;
        RECT 4.400 693.240 1558.640 694.640 ;
        RECT 4.000 689.200 1558.640 693.240 ;
        RECT 4.400 687.800 1558.640 689.200 ;
        RECT 4.000 683.760 1558.640 687.800 ;
        RECT 4.400 682.360 1558.640 683.760 ;
        RECT 4.000 678.320 1558.640 682.360 ;
        RECT 4.400 676.920 1558.640 678.320 ;
        RECT 4.000 672.880 1558.640 676.920 ;
        RECT 4.400 671.480 1558.640 672.880 ;
        RECT 4.000 667.440 1558.640 671.480 ;
        RECT 4.400 666.040 1558.640 667.440 ;
        RECT 4.000 662.000 1558.640 666.040 ;
        RECT 4.400 660.600 1558.640 662.000 ;
        RECT 4.000 656.560 1558.640 660.600 ;
        RECT 4.400 655.160 1558.640 656.560 ;
        RECT 4.000 651.120 1558.640 655.160 ;
        RECT 4.400 649.720 1558.640 651.120 ;
        RECT 4.000 645.680 1558.640 649.720 ;
        RECT 4.400 644.280 1558.640 645.680 ;
        RECT 4.000 640.920 1558.640 644.280 ;
        RECT 4.400 639.520 1558.640 640.920 ;
        RECT 4.000 635.480 1558.640 639.520 ;
        RECT 4.400 634.080 1558.640 635.480 ;
        RECT 4.000 630.040 1558.640 634.080 ;
        RECT 4.400 628.640 1558.640 630.040 ;
        RECT 4.000 624.600 1558.640 628.640 ;
        RECT 4.400 623.200 1558.640 624.600 ;
        RECT 4.000 619.160 1558.640 623.200 ;
        RECT 4.400 617.760 1558.640 619.160 ;
        RECT 4.000 613.720 1558.640 617.760 ;
        RECT 4.400 612.320 1558.640 613.720 ;
        RECT 4.000 608.280 1558.640 612.320 ;
        RECT 4.400 606.880 1558.640 608.280 ;
        RECT 4.000 602.840 1558.640 606.880 ;
        RECT 4.400 601.440 1558.640 602.840 ;
        RECT 4.000 597.400 1558.640 601.440 ;
        RECT 4.400 596.000 1558.640 597.400 ;
        RECT 4.000 591.960 1558.640 596.000 ;
        RECT 4.400 590.560 1558.640 591.960 ;
        RECT 4.000 586.520 1558.640 590.560 ;
        RECT 4.400 585.120 1558.640 586.520 ;
        RECT 4.000 581.080 1558.640 585.120 ;
        RECT 4.400 579.680 1558.640 581.080 ;
        RECT 4.000 575.640 1558.640 579.680 ;
        RECT 4.400 574.240 1558.640 575.640 ;
        RECT 4.000 570.200 1558.640 574.240 ;
        RECT 4.400 568.800 1558.640 570.200 ;
        RECT 4.000 564.760 1558.640 568.800 ;
        RECT 4.400 563.360 1558.640 564.760 ;
        RECT 4.000 559.320 1558.640 563.360 ;
        RECT 4.400 557.920 1558.640 559.320 ;
        RECT 4.000 553.880 1558.640 557.920 ;
        RECT 4.400 552.480 1558.640 553.880 ;
        RECT 4.000 548.440 1558.640 552.480 ;
        RECT 4.400 547.040 1558.640 548.440 ;
        RECT 4.000 543.000 1558.640 547.040 ;
        RECT 4.400 541.600 1558.640 543.000 ;
        RECT 4.000 537.560 1558.640 541.600 ;
        RECT 4.400 536.160 1558.640 537.560 ;
        RECT 4.000 532.800 1558.640 536.160 ;
        RECT 4.400 531.400 1558.640 532.800 ;
        RECT 4.000 527.360 1558.640 531.400 ;
        RECT 4.400 525.960 1558.640 527.360 ;
        RECT 4.000 521.920 1558.640 525.960 ;
        RECT 4.400 520.520 1558.640 521.920 ;
        RECT 4.000 516.480 1558.640 520.520 ;
        RECT 4.400 515.080 1558.640 516.480 ;
        RECT 4.000 511.040 1558.640 515.080 ;
        RECT 4.400 509.640 1558.640 511.040 ;
        RECT 4.000 505.600 1558.640 509.640 ;
        RECT 4.400 504.200 1558.640 505.600 ;
        RECT 4.000 500.160 1558.640 504.200 ;
        RECT 4.400 498.760 1558.640 500.160 ;
        RECT 4.000 494.720 1558.640 498.760 ;
        RECT 4.400 493.320 1558.640 494.720 ;
        RECT 4.000 489.280 1558.640 493.320 ;
        RECT 4.400 487.880 1558.640 489.280 ;
        RECT 4.000 483.840 1558.640 487.880 ;
        RECT 4.400 482.440 1558.640 483.840 ;
        RECT 4.000 478.400 1558.640 482.440 ;
        RECT 4.400 477.000 1558.640 478.400 ;
        RECT 4.000 472.960 1558.640 477.000 ;
        RECT 4.400 471.560 1558.640 472.960 ;
        RECT 4.000 467.520 1558.640 471.560 ;
        RECT 4.400 466.120 1558.640 467.520 ;
        RECT 4.000 462.080 1558.640 466.120 ;
        RECT 4.400 460.680 1558.640 462.080 ;
        RECT 4.000 456.640 1558.640 460.680 ;
        RECT 4.400 455.240 1558.640 456.640 ;
        RECT 4.000 451.200 1558.640 455.240 ;
        RECT 4.400 449.800 1558.640 451.200 ;
        RECT 4.000 445.760 1558.640 449.800 ;
        RECT 4.400 444.360 1558.640 445.760 ;
        RECT 4.000 440.320 1558.640 444.360 ;
        RECT 4.400 438.920 1558.640 440.320 ;
        RECT 4.000 434.880 1558.640 438.920 ;
        RECT 4.400 433.480 1558.640 434.880 ;
        RECT 4.000 429.440 1558.640 433.480 ;
        RECT 4.400 428.040 1558.640 429.440 ;
        RECT 4.000 424.680 1558.640 428.040 ;
        RECT 4.400 423.280 1558.640 424.680 ;
        RECT 4.000 419.240 1558.640 423.280 ;
        RECT 4.400 417.840 1558.640 419.240 ;
        RECT 4.000 413.800 1558.640 417.840 ;
        RECT 4.400 412.400 1558.640 413.800 ;
        RECT 4.000 408.360 1558.640 412.400 ;
        RECT 4.400 406.960 1558.640 408.360 ;
        RECT 4.000 402.920 1558.640 406.960 ;
        RECT 4.400 401.520 1558.640 402.920 ;
        RECT 4.000 397.480 1558.640 401.520 ;
        RECT 4.400 396.080 1558.640 397.480 ;
        RECT 4.000 392.040 1558.640 396.080 ;
        RECT 4.400 390.640 1558.640 392.040 ;
        RECT 4.000 386.600 1558.640 390.640 ;
        RECT 4.400 385.200 1558.640 386.600 ;
        RECT 4.000 381.160 1558.640 385.200 ;
        RECT 4.400 379.760 1558.640 381.160 ;
        RECT 4.000 375.720 1558.640 379.760 ;
        RECT 4.400 374.320 1558.640 375.720 ;
        RECT 4.000 370.280 1558.640 374.320 ;
        RECT 4.400 368.880 1558.640 370.280 ;
        RECT 4.000 364.840 1558.640 368.880 ;
        RECT 4.400 363.440 1558.640 364.840 ;
        RECT 4.000 359.400 1558.640 363.440 ;
        RECT 4.400 358.000 1558.640 359.400 ;
        RECT 4.000 353.960 1558.640 358.000 ;
        RECT 4.400 352.560 1558.640 353.960 ;
        RECT 4.000 348.520 1558.640 352.560 ;
        RECT 4.400 347.120 1558.640 348.520 ;
        RECT 4.000 343.080 1558.640 347.120 ;
        RECT 4.400 341.680 1558.640 343.080 ;
        RECT 4.000 337.640 1558.640 341.680 ;
        RECT 4.400 336.240 1558.640 337.640 ;
        RECT 4.000 332.200 1558.640 336.240 ;
        RECT 4.400 330.800 1558.640 332.200 ;
        RECT 4.000 326.760 1558.640 330.800 ;
        RECT 4.400 325.360 1558.640 326.760 ;
        RECT 4.000 322.000 1558.640 325.360 ;
        RECT 4.400 320.600 1558.640 322.000 ;
        RECT 4.000 316.560 1558.640 320.600 ;
        RECT 4.400 315.160 1558.640 316.560 ;
        RECT 4.000 311.120 1558.640 315.160 ;
        RECT 4.400 309.720 1558.640 311.120 ;
        RECT 4.000 305.680 1558.640 309.720 ;
        RECT 4.400 304.280 1558.640 305.680 ;
        RECT 4.000 300.240 1558.640 304.280 ;
        RECT 4.400 298.840 1558.640 300.240 ;
        RECT 4.000 294.800 1558.640 298.840 ;
        RECT 4.400 293.400 1558.640 294.800 ;
        RECT 4.000 289.360 1558.640 293.400 ;
        RECT 4.400 287.960 1558.640 289.360 ;
        RECT 4.000 283.920 1558.640 287.960 ;
        RECT 4.400 282.520 1558.640 283.920 ;
        RECT 4.000 278.480 1558.640 282.520 ;
        RECT 4.400 277.080 1558.640 278.480 ;
        RECT 4.000 273.040 1558.640 277.080 ;
        RECT 4.400 271.640 1558.640 273.040 ;
        RECT 4.000 267.600 1558.640 271.640 ;
        RECT 4.400 266.200 1558.640 267.600 ;
        RECT 4.000 262.160 1558.640 266.200 ;
        RECT 4.400 260.760 1558.640 262.160 ;
        RECT 4.000 256.720 1558.640 260.760 ;
        RECT 4.400 255.320 1558.640 256.720 ;
        RECT 4.000 251.280 1558.640 255.320 ;
        RECT 4.400 249.880 1558.640 251.280 ;
        RECT 4.000 245.840 1558.640 249.880 ;
        RECT 4.400 244.440 1558.640 245.840 ;
        RECT 4.000 240.400 1558.640 244.440 ;
        RECT 4.400 239.000 1558.640 240.400 ;
        RECT 4.000 234.960 1558.640 239.000 ;
        RECT 4.400 233.560 1558.640 234.960 ;
        RECT 4.000 229.520 1558.640 233.560 ;
        RECT 4.400 228.120 1558.640 229.520 ;
        RECT 4.000 224.080 1558.640 228.120 ;
        RECT 4.400 222.680 1558.640 224.080 ;
        RECT 4.000 218.640 1558.640 222.680 ;
        RECT 4.400 217.240 1558.640 218.640 ;
        RECT 4.000 213.880 1558.640 217.240 ;
        RECT 4.400 212.480 1558.640 213.880 ;
        RECT 4.000 208.440 1558.640 212.480 ;
        RECT 4.400 207.040 1558.640 208.440 ;
        RECT 4.000 203.000 1558.640 207.040 ;
        RECT 4.400 201.600 1558.640 203.000 ;
        RECT 4.000 197.560 1558.640 201.600 ;
        RECT 4.400 196.160 1558.640 197.560 ;
        RECT 4.000 192.120 1558.640 196.160 ;
        RECT 4.400 190.720 1558.640 192.120 ;
        RECT 4.000 186.680 1558.640 190.720 ;
        RECT 4.400 185.280 1558.640 186.680 ;
        RECT 4.000 181.240 1558.640 185.280 ;
        RECT 4.400 179.840 1558.640 181.240 ;
        RECT 4.000 175.800 1558.640 179.840 ;
        RECT 4.400 174.400 1558.640 175.800 ;
        RECT 4.000 170.360 1558.640 174.400 ;
        RECT 4.400 168.960 1558.640 170.360 ;
        RECT 4.000 164.920 1558.640 168.960 ;
        RECT 4.400 163.520 1558.640 164.920 ;
        RECT 4.000 159.480 1558.640 163.520 ;
        RECT 4.400 158.080 1558.640 159.480 ;
        RECT 4.000 154.040 1558.640 158.080 ;
        RECT 4.400 152.640 1558.640 154.040 ;
        RECT 4.000 148.600 1558.640 152.640 ;
        RECT 4.400 147.200 1558.640 148.600 ;
        RECT 4.000 143.160 1558.640 147.200 ;
        RECT 4.400 141.760 1558.640 143.160 ;
        RECT 4.000 137.720 1558.640 141.760 ;
        RECT 4.400 136.320 1558.640 137.720 ;
        RECT 4.000 132.280 1558.640 136.320 ;
        RECT 4.400 130.880 1558.640 132.280 ;
        RECT 4.000 126.840 1558.640 130.880 ;
        RECT 4.400 125.440 1558.640 126.840 ;
        RECT 4.000 121.400 1558.640 125.440 ;
        RECT 4.400 120.000 1558.640 121.400 ;
        RECT 4.000 115.960 1558.640 120.000 ;
        RECT 4.400 114.560 1558.640 115.960 ;
        RECT 4.000 110.520 1558.640 114.560 ;
        RECT 4.400 109.120 1558.640 110.520 ;
        RECT 4.000 105.760 1558.640 109.120 ;
        RECT 4.400 104.360 1558.640 105.760 ;
        RECT 4.000 100.320 1558.640 104.360 ;
        RECT 4.400 98.920 1558.640 100.320 ;
        RECT 4.000 94.880 1558.640 98.920 ;
        RECT 4.400 93.480 1558.640 94.880 ;
        RECT 4.000 89.440 1558.640 93.480 ;
        RECT 4.400 88.040 1558.640 89.440 ;
        RECT 4.000 84.000 1558.640 88.040 ;
        RECT 4.400 82.600 1558.640 84.000 ;
        RECT 4.000 78.560 1558.640 82.600 ;
        RECT 4.400 77.160 1558.640 78.560 ;
        RECT 4.000 73.120 1558.640 77.160 ;
        RECT 4.400 71.720 1558.640 73.120 ;
        RECT 4.000 67.680 1558.640 71.720 ;
        RECT 4.400 66.280 1558.640 67.680 ;
        RECT 4.000 62.240 1558.640 66.280 ;
        RECT 4.400 60.840 1558.640 62.240 ;
        RECT 4.000 56.800 1558.640 60.840 ;
        RECT 4.400 55.400 1558.640 56.800 ;
        RECT 4.000 51.360 1558.640 55.400 ;
        RECT 4.400 49.960 1558.640 51.360 ;
        RECT 4.000 45.920 1558.640 49.960 ;
        RECT 4.400 44.520 1558.640 45.920 ;
        RECT 4.000 40.480 1558.640 44.520 ;
        RECT 4.400 39.080 1558.640 40.480 ;
        RECT 4.000 35.040 1558.640 39.080 ;
        RECT 4.400 33.640 1558.640 35.040 ;
        RECT 4.000 29.600 1558.640 33.640 ;
        RECT 4.400 28.200 1558.640 29.600 ;
        RECT 4.000 24.160 1558.640 28.200 ;
        RECT 4.400 22.760 1558.640 24.160 ;
        RECT 4.000 18.720 1558.640 22.760 ;
        RECT 4.400 17.320 1558.640 18.720 ;
        RECT 4.000 13.280 1558.640 17.320 ;
        RECT 4.400 11.880 1558.640 13.280 ;
        RECT 4.000 7.840 1558.640 11.880 ;
        RECT 4.400 6.440 1558.640 7.840 ;
        RECT 4.000 3.080 1558.640 6.440 ;
        RECT 4.400 2.215 1558.640 3.080 ;
      LAYER met4 ;
        RECT 4.895 12.415 20.640 1587.625 ;
        RECT 23.040 12.415 97.440 1587.625 ;
        RECT 99.840 12.415 174.240 1587.625 ;
        RECT 176.640 12.415 251.040 1587.625 ;
        RECT 253.440 12.415 327.840 1587.625 ;
        RECT 330.240 12.415 404.640 1587.625 ;
        RECT 407.040 12.415 481.440 1587.625 ;
        RECT 483.840 12.415 558.240 1587.625 ;
        RECT 560.640 12.415 635.040 1587.625 ;
        RECT 637.440 12.415 711.840 1587.625 ;
        RECT 714.240 12.415 788.640 1587.625 ;
        RECT 791.040 12.415 844.265 1587.625 ;
  END
END c0_system
END LIBRARY


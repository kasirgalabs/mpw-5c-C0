VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO c0_system
  CLASS BLOCK ;
  FOREIGN c0_system ;
  ORIGIN 0.000 0.000 ;
  SIZE 1300.000 BY 1300.000 ;
  PIN bb_addr0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 581.440 4.000 582.040 ;
    END
  END bb_addr0[0]
  PIN bb_addr0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 818.760 4.000 819.360 ;
    END
  END bb_addr0[10]
  PIN bb_addr0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 840.520 4.000 841.120 ;
    END
  END bb_addr0[11]
  PIN bb_addr0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 862.960 4.000 863.560 ;
    END
  END bb_addr0[12]
  PIN bb_addr0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 884.720 4.000 885.320 ;
    END
  END bb_addr0[13]
  PIN bb_addr0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 906.480 4.000 907.080 ;
    END
  END bb_addr0[14]
  PIN bb_addr0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 928.240 4.000 928.840 ;
    END
  END bb_addr0[15]
  PIN bb_addr0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 950.680 4.000 951.280 ;
    END
  END bb_addr0[16]
  PIN bb_addr0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 972.440 4.000 973.040 ;
    END
  END bb_addr0[17]
  PIN bb_addr0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 994.200 4.000 994.800 ;
    END
  END bb_addr0[18]
  PIN bb_addr0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1016.640 4.000 1017.240 ;
    END
  END bb_addr0[19]
  PIN bb_addr0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 607.960 4.000 608.560 ;
    END
  END bb_addr0[1]
  PIN bb_addr0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1038.400 4.000 1039.000 ;
    END
  END bb_addr0[20]
  PIN bb_addr0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1060.160 4.000 1060.760 ;
    END
  END bb_addr0[21]
  PIN bb_addr0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1082.600 4.000 1083.200 ;
    END
  END bb_addr0[22]
  PIN bb_addr0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1104.360 4.000 1104.960 ;
    END
  END bb_addr0[23]
  PIN bb_addr0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1126.120 4.000 1126.720 ;
    END
  END bb_addr0[24]
  PIN bb_addr0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1147.880 4.000 1148.480 ;
    END
  END bb_addr0[25]
  PIN bb_addr0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1170.320 4.000 1170.920 ;
    END
  END bb_addr0[26]
  PIN bb_addr0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1192.080 4.000 1192.680 ;
    END
  END bb_addr0[27]
  PIN bb_addr0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1213.840 4.000 1214.440 ;
    END
  END bb_addr0[28]
  PIN bb_addr0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1236.280 4.000 1236.880 ;
    END
  END bb_addr0[29]
  PIN bb_addr0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 634.480 4.000 635.080 ;
    END
  END bb_addr0[2]
  PIN bb_addr0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1258.040 4.000 1258.640 ;
    END
  END bb_addr0[30]
  PIN bb_addr0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1279.800 4.000 1280.400 ;
    END
  END bb_addr0[31]
  PIN bb_addr0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 660.320 4.000 660.920 ;
    END
  END bb_addr0[3]
  PIN bb_addr0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 686.840 4.000 687.440 ;
    END
  END bb_addr0[4]
  PIN bb_addr0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 708.600 4.000 709.200 ;
    END
  END bb_addr0[5]
  PIN bb_addr0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 731.040 4.000 731.640 ;
    END
  END bb_addr0[6]
  PIN bb_addr0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 752.800 4.000 753.400 ;
    END
  END bb_addr0[7]
  PIN bb_addr0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 774.560 4.000 775.160 ;
    END
  END bb_addr0[8]
  PIN bb_addr0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 797.000 4.000 797.600 ;
    END
  END bb_addr0[9]
  PIN bb_addr1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 586.200 4.000 586.800 ;
    END
  END bb_addr1[0]
  PIN bb_addr1[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 822.840 4.000 823.440 ;
    END
  END bb_addr1[10]
  PIN bb_addr1[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 845.280 4.000 845.880 ;
    END
  END bb_addr1[11]
  PIN bb_addr1[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 867.040 4.000 867.640 ;
    END
  END bb_addr1[12]
  PIN bb_addr1[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 888.800 4.000 889.400 ;
    END
  END bb_addr1[13]
  PIN bb_addr1[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 911.240 4.000 911.840 ;
    END
  END bb_addr1[14]
  PIN bb_addr1[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 933.000 4.000 933.600 ;
    END
  END bb_addr1[15]
  PIN bb_addr1[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 954.760 4.000 955.360 ;
    END
  END bb_addr1[16]
  PIN bb_addr1[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 977.200 4.000 977.800 ;
    END
  END bb_addr1[17]
  PIN bb_addr1[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 998.960 4.000 999.560 ;
    END
  END bb_addr1[18]
  PIN bb_addr1[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1020.720 4.000 1021.320 ;
    END
  END bb_addr1[19]
  PIN bb_addr1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 612.040 4.000 612.640 ;
    END
  END bb_addr1[1]
  PIN bb_addr1[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1042.480 4.000 1043.080 ;
    END
  END bb_addr1[20]
  PIN bb_addr1[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1064.920 4.000 1065.520 ;
    END
  END bb_addr1[21]
  PIN bb_addr1[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1086.680 4.000 1087.280 ;
    END
  END bb_addr1[22]
  PIN bb_addr1[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1108.440 4.000 1109.040 ;
    END
  END bb_addr1[23]
  PIN bb_addr1[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1130.880 4.000 1131.480 ;
    END
  END bb_addr1[24]
  PIN bb_addr1[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1152.640 4.000 1153.240 ;
    END
  END bb_addr1[25]
  PIN bb_addr1[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1174.400 4.000 1175.000 ;
    END
  END bb_addr1[26]
  PIN bb_addr1[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1196.160 4.000 1196.760 ;
    END
  END bb_addr1[27]
  PIN bb_addr1[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1218.600 4.000 1219.200 ;
    END
  END bb_addr1[28]
  PIN bb_addr1[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1240.360 4.000 1240.960 ;
    END
  END bb_addr1[29]
  PIN bb_addr1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 638.560 4.000 639.160 ;
    END
  END bb_addr1[2]
  PIN bb_addr1[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1262.120 4.000 1262.720 ;
    END
  END bb_addr1[30]
  PIN bb_addr1[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1284.560 4.000 1285.160 ;
    END
  END bb_addr1[31]
  PIN bb_addr1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 665.080 4.000 665.680 ;
    END
  END bb_addr1[3]
  PIN bb_addr1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 691.600 4.000 692.200 ;
    END
  END bb_addr1[4]
  PIN bb_addr1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 713.360 4.000 713.960 ;
    END
  END bb_addr1[5]
  PIN bb_addr1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 735.120 4.000 735.720 ;
    END
  END bb_addr1[6]
  PIN bb_addr1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 757.560 4.000 758.160 ;
    END
  END bb_addr1[7]
  PIN bb_addr1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 779.320 4.000 779.920 ;
    END
  END bb_addr1[8]
  PIN bb_addr1[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 801.080 4.000 801.680 ;
    END
  END bb_addr1[9]
  PIN bb_csb0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 568.520 4.000 569.120 ;
    END
  END bb_csb0
  PIN bb_csb1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 572.600 4.000 573.200 ;
    END
  END bb_csb1
  PIN bb_din0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 590.280 4.000 590.880 ;
    END
  END bb_din0[0]
  PIN bb_din0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 827.600 4.000 828.200 ;
    END
  END bb_din0[10]
  PIN bb_din0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 849.360 4.000 849.960 ;
    END
  END bb_din0[11]
  PIN bb_din0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 871.120 4.000 871.720 ;
    END
  END bb_din0[12]
  PIN bb_din0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 893.560 4.000 894.160 ;
    END
  END bb_din0[13]
  PIN bb_din0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 915.320 4.000 915.920 ;
    END
  END bb_din0[14]
  PIN bb_din0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 937.080 4.000 937.680 ;
    END
  END bb_din0[15]
  PIN bb_din0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 959.520 4.000 960.120 ;
    END
  END bb_din0[16]
  PIN bb_din0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 981.280 4.000 981.880 ;
    END
  END bb_din0[17]
  PIN bb_din0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1003.040 4.000 1003.640 ;
    END
  END bb_din0[18]
  PIN bb_din0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1025.480 4.000 1026.080 ;
    END
  END bb_din0[19]
  PIN bb_din0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 616.800 4.000 617.400 ;
    END
  END bb_din0[1]
  PIN bb_din0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1047.240 4.000 1047.840 ;
    END
  END bb_din0[20]
  PIN bb_din0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1069.000 4.000 1069.600 ;
    END
  END bb_din0[21]
  PIN bb_din0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1090.760 4.000 1091.360 ;
    END
  END bb_din0[22]
  PIN bb_din0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1113.200 4.000 1113.800 ;
    END
  END bb_din0[23]
  PIN bb_din0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1134.960 4.000 1135.560 ;
    END
  END bb_din0[24]
  PIN bb_din0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1156.720 4.000 1157.320 ;
    END
  END bb_din0[25]
  PIN bb_din0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1179.160 4.000 1179.760 ;
    END
  END bb_din0[26]
  PIN bb_din0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1200.920 4.000 1201.520 ;
    END
  END bb_din0[27]
  PIN bb_din0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1222.680 4.000 1223.280 ;
    END
  END bb_din0[28]
  PIN bb_din0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1245.120 4.000 1245.720 ;
    END
  END bb_din0[29]
  PIN bb_din0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 643.320 4.000 643.920 ;
    END
  END bb_din0[2]
  PIN bb_din0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1266.880 4.000 1267.480 ;
    END
  END bb_din0[30]
  PIN bb_din0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1288.640 4.000 1289.240 ;
    END
  END bb_din0[31]
  PIN bb_din0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 669.160 4.000 669.760 ;
    END
  END bb_din0[3]
  PIN bb_din0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 695.680 4.000 696.280 ;
    END
  END bb_din0[4]
  PIN bb_din0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 717.440 4.000 718.040 ;
    END
  END bb_din0[5]
  PIN bb_din0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 739.880 4.000 740.480 ;
    END
  END bb_din0[6]
  PIN bb_din0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 761.640 4.000 762.240 ;
    END
  END bb_din0[7]
  PIN bb_din0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 783.400 4.000 784.000 ;
    END
  END bb_din0[8]
  PIN bb_din0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 805.840 4.000 806.440 ;
    END
  END bb_din0[9]
  PIN bb_dout0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 595.040 4.000 595.640 ;
    END
  END bb_dout0[0]
  PIN bb_dout0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 831.680 4.000 832.280 ;
    END
  END bb_dout0[10]
  PIN bb_dout0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 854.120 4.000 854.720 ;
    END
  END bb_dout0[11]
  PIN bb_dout0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 875.880 4.000 876.480 ;
    END
  END bb_dout0[12]
  PIN bb_dout0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 897.640 4.000 898.240 ;
    END
  END bb_dout0[13]
  PIN bb_dout0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 920.080 4.000 920.680 ;
    END
  END bb_dout0[14]
  PIN bb_dout0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 941.840 4.000 942.440 ;
    END
  END bb_dout0[15]
  PIN bb_dout0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 963.600 4.000 964.200 ;
    END
  END bb_dout0[16]
  PIN bb_dout0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 985.360 4.000 985.960 ;
    END
  END bb_dout0[17]
  PIN bb_dout0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1007.800 4.000 1008.400 ;
    END
  END bb_dout0[18]
  PIN bb_dout0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1029.560 4.000 1030.160 ;
    END
  END bb_dout0[19]
  PIN bb_dout0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 620.880 4.000 621.480 ;
    END
  END bb_dout0[1]
  PIN bb_dout0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1051.320 4.000 1051.920 ;
    END
  END bb_dout0[20]
  PIN bb_dout0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1073.760 4.000 1074.360 ;
    END
  END bb_dout0[21]
  PIN bb_dout0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1095.520 4.000 1096.120 ;
    END
  END bb_dout0[22]
  PIN bb_dout0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1117.280 4.000 1117.880 ;
    END
  END bb_dout0[23]
  PIN bb_dout0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1139.720 4.000 1140.320 ;
    END
  END bb_dout0[24]
  PIN bb_dout0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1161.480 4.000 1162.080 ;
    END
  END bb_dout0[25]
  PIN bb_dout0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1183.240 4.000 1183.840 ;
    END
  END bb_dout0[26]
  PIN bb_dout0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1205.000 4.000 1205.600 ;
    END
  END bb_dout0[27]
  PIN bb_dout0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1227.440 4.000 1228.040 ;
    END
  END bb_dout0[28]
  PIN bb_dout0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1249.200 4.000 1249.800 ;
    END
  END bb_dout0[29]
  PIN bb_dout0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 647.400 4.000 648.000 ;
    END
  END bb_dout0[2]
  PIN bb_dout0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1270.960 4.000 1271.560 ;
    END
  END bb_dout0[30]
  PIN bb_dout0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1293.400 4.000 1294.000 ;
    END
  END bb_dout0[31]
  PIN bb_dout0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 673.920 4.000 674.520 ;
    END
  END bb_dout0[3]
  PIN bb_dout0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 700.440 4.000 701.040 ;
    END
  END bb_dout0[4]
  PIN bb_dout0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 722.200 4.000 722.800 ;
    END
  END bb_dout0[5]
  PIN bb_dout0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 743.960 4.000 744.560 ;
    END
  END bb_dout0[6]
  PIN bb_dout0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 765.720 4.000 766.320 ;
    END
  END bb_dout0[7]
  PIN bb_dout0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 788.160 4.000 788.760 ;
    END
  END bb_dout0[8]
  PIN bb_dout0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 809.920 4.000 810.520 ;
    END
  END bb_dout0[9]
  PIN bb_dout1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 599.120 4.000 599.720 ;
    END
  END bb_dout1[0]
  PIN bb_dout1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 836.440 4.000 837.040 ;
    END
  END bb_dout1[10]
  PIN bb_dout1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 858.200 4.000 858.800 ;
    END
  END bb_dout1[11]
  PIN bb_dout1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 879.960 4.000 880.560 ;
    END
  END bb_dout1[12]
  PIN bb_dout1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 902.400 4.000 903.000 ;
    END
  END bb_dout1[13]
  PIN bb_dout1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 924.160 4.000 924.760 ;
    END
  END bb_dout1[14]
  PIN bb_dout1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 945.920 4.000 946.520 ;
    END
  END bb_dout1[15]
  PIN bb_dout1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 968.360 4.000 968.960 ;
    END
  END bb_dout1[16]
  PIN bb_dout1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 990.120 4.000 990.720 ;
    END
  END bb_dout1[17]
  PIN bb_dout1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1011.880 4.000 1012.480 ;
    END
  END bb_dout1[18]
  PIN bb_dout1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1033.640 4.000 1034.240 ;
    END
  END bb_dout1[19]
  PIN bb_dout1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 625.640 4.000 626.240 ;
    END
  END bb_dout1[1]
  PIN bb_dout1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1056.080 4.000 1056.680 ;
    END
  END bb_dout1[20]
  PIN bb_dout1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1077.840 4.000 1078.440 ;
    END
  END bb_dout1[21]
  PIN bb_dout1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1099.600 4.000 1100.200 ;
    END
  END bb_dout1[22]
  PIN bb_dout1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1122.040 4.000 1122.640 ;
    END
  END bb_dout1[23]
  PIN bb_dout1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1143.800 4.000 1144.400 ;
    END
  END bb_dout1[24]
  PIN bb_dout1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1165.560 4.000 1166.160 ;
    END
  END bb_dout1[25]
  PIN bb_dout1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1188.000 4.000 1188.600 ;
    END
  END bb_dout1[26]
  PIN bb_dout1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1209.760 4.000 1210.360 ;
    END
  END bb_dout1[27]
  PIN bb_dout1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1231.520 4.000 1232.120 ;
    END
  END bb_dout1[28]
  PIN bb_dout1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1253.280 4.000 1253.880 ;
    END
  END bb_dout1[29]
  PIN bb_dout1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 652.160 4.000 652.760 ;
    END
  END bb_dout1[2]
  PIN bb_dout1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1275.720 4.000 1276.320 ;
    END
  END bb_dout1[30]
  PIN bb_dout1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1297.480 4.000 1298.080 ;
    END
  END bb_dout1[31]
  PIN bb_dout1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 678.000 4.000 678.600 ;
    END
  END bb_dout1[3]
  PIN bb_dout1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 704.520 4.000 705.120 ;
    END
  END bb_dout1[4]
  PIN bb_dout1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 726.280 4.000 726.880 ;
    END
  END bb_dout1[5]
  PIN bb_dout1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 748.720 4.000 749.320 ;
    END
  END bb_dout1[6]
  PIN bb_dout1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 770.480 4.000 771.080 ;
    END
  END bb_dout1[7]
  PIN bb_dout1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 792.240 4.000 792.840 ;
    END
  END bb_dout1[8]
  PIN bb_dout1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 814.680 4.000 815.280 ;
    END
  END bb_dout1[9]
  PIN bb_web0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 577.360 4.000 577.960 ;
    END
  END bb_web0
  PIN bb_wmask0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 603.200 4.000 603.800 ;
    END
  END bb_wmask0[0]
  PIN bb_wmask0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 629.720 4.000 630.320 ;
    END
  END bb_wmask0[1]
  PIN bb_wmask0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 656.240 4.000 656.840 ;
    END
  END bb_wmask0[2]
  PIN bb_wmask0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 682.760 4.000 683.360 ;
    END
  END bb_wmask0[3]
  PIN clk_g
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.370 0.000 8.650 4.000 ;
    END
  END clk_g
  PIN io_gecerli
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 4.000 ;
    END
  END io_gecerli
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.850 0.000 95.130 4.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.690 0.000 441.970 4.000 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 476.190 0.000 476.470 4.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 510.690 0.000 510.970 4.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 545.650 0.000 545.930 4.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 580.150 0.000 580.430 4.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 614.650 0.000 614.930 4.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 649.610 0.000 649.890 4.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 684.110 0.000 684.390 4.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 718.610 0.000 718.890 4.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 753.570 0.000 753.850 4.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.350 0.000 129.630 4.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 788.070 0.000 788.350 4.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 822.570 0.000 822.850 4.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 857.530 0.000 857.810 4.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 892.030 0.000 892.310 4.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 926.990 0.000 927.270 4.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 961.490 0.000 961.770 4.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 995.990 0.000 996.270 4.000 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1030.950 0.000 1031.230 4.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1065.450 0.000 1065.730 4.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1099.950 0.000 1100.230 4.000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 0.000 164.590 4.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1134.910 0.000 1135.190 4.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1169.410 0.000 1169.690 4.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1203.910 0.000 1204.190 4.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1221.390 0.000 1221.670 4.000 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1238.870 0.000 1239.150 4.000 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1255.890 0.000 1256.170 4.000 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1273.370 0.000 1273.650 4.000 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1290.850 0.000 1291.130 4.000 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.810 0.000 199.090 4.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.310 0.000 233.590 4.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.270 0.000 268.550 4.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.770 0.000 303.050 4.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 337.270 0.000 337.550 4.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 372.230 0.000 372.510 4.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 406.730 0.000 407.010 4.000 ;
    END
  END io_oeb[9]
  PIN io_ps[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.330 0.000 112.610 4.000 ;
    END
  END io_ps[0]
  PIN io_ps[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 458.710 0.000 458.990 4.000 ;
    END
  END io_ps[10]
  PIN io_ps[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 493.670 0.000 493.950 4.000 ;
    END
  END io_ps[11]
  PIN io_ps[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.170 0.000 528.450 4.000 ;
    END
  END io_ps[12]
  PIN io_ps[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 562.670 0.000 562.950 4.000 ;
    END
  END io_ps[13]
  PIN io_ps[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 597.630 0.000 597.910 4.000 ;
    END
  END io_ps[14]
  PIN io_ps[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 632.130 0.000 632.410 4.000 ;
    END
  END io_ps[15]
  PIN io_ps[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 666.630 0.000 666.910 4.000 ;
    END
  END io_ps[16]
  PIN io_ps[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 701.590 0.000 701.870 4.000 ;
    END
  END io_ps[17]
  PIN io_ps[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 736.090 0.000 736.370 4.000 ;
    END
  END io_ps[18]
  PIN io_ps[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 770.590 0.000 770.870 4.000 ;
    END
  END io_ps[19]
  PIN io_ps[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.830 0.000 147.110 4.000 ;
    END
  END io_ps[1]
  PIN io_ps[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 805.550 0.000 805.830 4.000 ;
    END
  END io_ps[20]
  PIN io_ps[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 840.050 0.000 840.330 4.000 ;
    END
  END io_ps[21]
  PIN io_ps[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 875.010 0.000 875.290 4.000 ;
    END
  END io_ps[22]
  PIN io_ps[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 909.510 0.000 909.790 4.000 ;
    END
  END io_ps[23]
  PIN io_ps[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 944.010 0.000 944.290 4.000 ;
    END
  END io_ps[24]
  PIN io_ps[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 978.970 0.000 979.250 4.000 ;
    END
  END io_ps[25]
  PIN io_ps[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1013.470 0.000 1013.750 4.000 ;
    END
  END io_ps[26]
  PIN io_ps[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1047.970 0.000 1048.250 4.000 ;
    END
  END io_ps[27]
  PIN io_ps[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1082.930 0.000 1083.210 4.000 ;
    END
  END io_ps[28]
  PIN io_ps[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1117.430 0.000 1117.710 4.000 ;
    END
  END io_ps[29]
  PIN io_ps[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.330 0.000 181.610 4.000 ;
    END
  END io_ps[2]
  PIN io_ps[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1151.930 0.000 1152.210 4.000 ;
    END
  END io_ps[30]
  PIN io_ps[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1186.890 0.000 1187.170 4.000 ;
    END
  END io_ps[31]
  PIN io_ps[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.290 0.000 216.570 4.000 ;
    END
  END io_ps[3]
  PIN io_ps[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.790 0.000 251.070 4.000 ;
    END
  END io_ps[4]
  PIN io_ps[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.290 0.000 285.570 4.000 ;
    END
  END io_ps[5]
  PIN io_ps[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 320.250 0.000 320.530 4.000 ;
    END
  END io_ps[6]
  PIN io_ps[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.750 0.000 355.030 4.000 ;
    END
  END io_ps[7]
  PIN io_ps[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.250 0.000 389.530 4.000 ;
    END
  END io_ps[8]
  PIN io_ps[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 424.210 0.000 424.490 4.000 ;
    END
  END io_ps[9]
  PIN rst_g
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.390 0.000 25.670 4.000 ;
    END
  END rst_g
  PIN rx
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.350 0.000 60.630 4.000 ;
    END
  END rx
  PIN tx
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.870 0.000 43.150 4.000 ;
    END
  END tx
  PIN vb_addr0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.000 4.000 15.600 ;
    END
  END vb_addr0[0]
  PIN vb_addr0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 252.320 4.000 252.920 ;
    END
  END vb_addr0[10]
  PIN vb_addr0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 274.080 4.000 274.680 ;
    END
  END vb_addr0[11]
  PIN vb_addr0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 295.840 4.000 296.440 ;
    END
  END vb_addr0[12]
  PIN vb_addr0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 41.520 4.000 42.120 ;
    END
  END vb_addr0[1]
  PIN vb_addr0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 67.360 4.000 67.960 ;
    END
  END vb_addr0[2]
  PIN vb_addr0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.880 4.000 94.480 ;
    END
  END vb_addr0[3]
  PIN vb_addr0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 120.400 4.000 121.000 ;
    END
  END vb_addr0[4]
  PIN vb_addr0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.160 4.000 142.760 ;
    END
  END vb_addr0[5]
  PIN vb_addr0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 164.600 4.000 165.200 ;
    END
  END vb_addr0[6]
  PIN vb_addr0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 186.360 4.000 186.960 ;
    END
  END vb_addr0[7]
  PIN vb_addr0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 208.120 4.000 208.720 ;
    END
  END vb_addr0[8]
  PIN vb_addr0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 229.880 4.000 230.480 ;
    END
  END vb_addr0[9]
  PIN vb_addr1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.080 4.000 19.680 ;
    END
  END vb_addr1[0]
  PIN vb_addr1[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 256.400 4.000 257.000 ;
    END
  END vb_addr1[10]
  PIN vb_addr1[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 278.160 4.000 278.760 ;
    END
  END vb_addr1[11]
  PIN vb_addr1[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 300.600 4.000 301.200 ;
    END
  END vb_addr1[12]
  PIN vb_addr1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 45.600 4.000 46.200 ;
    END
  END vb_addr1[1]
  PIN vb_addr1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.120 4.000 72.720 ;
    END
  END vb_addr1[2]
  PIN vb_addr1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 98.640 4.000 99.240 ;
    END
  END vb_addr1[3]
  PIN vb_addr1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 124.480 4.000 125.080 ;
    END
  END vb_addr1[4]
  PIN vb_addr1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.920 4.000 147.520 ;
    END
  END vb_addr1[5]
  PIN vb_addr1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.680 4.000 169.280 ;
    END
  END vb_addr1[6]
  PIN vb_addr1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 190.440 4.000 191.040 ;
    END
  END vb_addr1[7]
  PIN vb_addr1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 212.880 4.000 213.480 ;
    END
  END vb_addr1[8]
  PIN vb_addr1[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 234.640 4.000 235.240 ;
    END
  END vb_addr1[9]
  PIN vb_csb0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.080 4.000 2.680 ;
    END
  END vb_csb0
  PIN vb_csb1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.160 4.000 6.760 ;
    END
  END vb_csb1
  PIN vb_din0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 4.000 24.440 ;
    END
  END vb_din0[0]
  PIN vb_din0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 261.160 4.000 261.760 ;
    END
  END vb_din0[10]
  PIN vb_din0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 282.920 4.000 283.520 ;
    END
  END vb_din0[11]
  PIN vb_din0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 304.680 4.000 305.280 ;
    END
  END vb_din0[12]
  PIN vb_din0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 318.280 4.000 318.880 ;
    END
  END vb_din0[13]
  PIN vb_din0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 331.200 4.000 331.800 ;
    END
  END vb_din0[14]
  PIN vb_din0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 344.120 4.000 344.720 ;
    END
  END vb_din0[15]
  PIN vb_din0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 357.720 4.000 358.320 ;
    END
  END vb_din0[16]
  PIN vb_din0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 370.640 4.000 371.240 ;
    END
  END vb_din0[17]
  PIN vb_din0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 383.560 4.000 384.160 ;
    END
  END vb_din0[18]
  PIN vb_din0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 397.160 4.000 397.760 ;
    END
  END vb_din0[19]
  PIN vb_din0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 50.360 4.000 50.960 ;
    END
  END vb_din0[1]
  PIN vb_din0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 410.080 4.000 410.680 ;
    END
  END vb_din0[20]
  PIN vb_din0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 423.680 4.000 424.280 ;
    END
  END vb_din0[21]
  PIN vb_din0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 436.600 4.000 437.200 ;
    END
  END vb_din0[22]
  PIN vb_din0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 449.520 4.000 450.120 ;
    END
  END vb_din0[23]
  PIN vb_din0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 463.120 4.000 463.720 ;
    END
  END vb_din0[24]
  PIN vb_din0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 476.040 4.000 476.640 ;
    END
  END vb_din0[25]
  PIN vb_din0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 489.640 4.000 490.240 ;
    END
  END vb_din0[26]
  PIN vb_din0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 502.560 4.000 503.160 ;
    END
  END vb_din0[27]
  PIN vb_din0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 515.480 4.000 516.080 ;
    END
  END vb_din0[28]
  PIN vb_din0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 529.080 4.000 529.680 ;
    END
  END vb_din0[29]
  PIN vb_din0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.200 4.000 76.800 ;
    END
  END vb_din0[2]
  PIN vb_din0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 542.000 4.000 542.600 ;
    END
  END vb_din0[30]
  PIN vb_din0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 554.920 4.000 555.520 ;
    END
  END vb_din0[31]
  PIN vb_din0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.720 4.000 103.320 ;
    END
  END vb_din0[3]
  PIN vb_din0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 4.000 129.840 ;
    END
  END vb_din0[4]
  PIN vb_din0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 151.000 4.000 151.600 ;
    END
  END vb_din0[5]
  PIN vb_din0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 172.760 4.000 173.360 ;
    END
  END vb_din0[6]
  PIN vb_din0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 195.200 4.000 195.800 ;
    END
  END vb_din0[7]
  PIN vb_din0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 216.960 4.000 217.560 ;
    END
  END vb_din0[8]
  PIN vb_din0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 238.720 4.000 239.320 ;
    END
  END vb_din0[9]
  PIN vb_dout0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.920 4.000 28.520 ;
    END
  END vb_dout0[0]
  PIN vb_dout0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 265.240 4.000 265.840 ;
    END
  END vb_dout0[10]
  PIN vb_dout0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 287.000 4.000 287.600 ;
    END
  END vb_dout0[11]
  PIN vb_dout0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 309.440 4.000 310.040 ;
    END
  END vb_dout0[12]
  PIN vb_dout0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 322.360 4.000 322.960 ;
    END
  END vb_dout0[13]
  PIN vb_dout0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 335.280 4.000 335.880 ;
    END
  END vb_dout0[14]
  PIN vb_dout0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 348.880 4.000 349.480 ;
    END
  END vb_dout0[15]
  PIN vb_dout0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 361.800 4.000 362.400 ;
    END
  END vb_dout0[16]
  PIN vb_dout0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 375.400 4.000 376.000 ;
    END
  END vb_dout0[17]
  PIN vb_dout0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 388.320 4.000 388.920 ;
    END
  END vb_dout0[18]
  PIN vb_dout0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 401.240 4.000 401.840 ;
    END
  END vb_dout0[19]
  PIN vb_dout0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END vb_dout0[1]
  PIN vb_dout0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 414.840 4.000 415.440 ;
    END
  END vb_dout0[20]
  PIN vb_dout0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 427.760 4.000 428.360 ;
    END
  END vb_dout0[21]
  PIN vb_dout0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 440.680 4.000 441.280 ;
    END
  END vb_dout0[22]
  PIN vb_dout0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 454.280 4.000 454.880 ;
    END
  END vb_dout0[23]
  PIN vb_dout0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 467.200 4.000 467.800 ;
    END
  END vb_dout0[24]
  PIN vb_dout0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 480.800 4.000 481.400 ;
    END
  END vb_dout0[25]
  PIN vb_dout0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 493.720 4.000 494.320 ;
    END
  END vb_dout0[26]
  PIN vb_dout0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 506.640 4.000 507.240 ;
    END
  END vb_dout0[27]
  PIN vb_dout0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 520.240 4.000 520.840 ;
    END
  END vb_dout0[28]
  PIN vb_dout0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 533.160 4.000 533.760 ;
    END
  END vb_dout0[29]
  PIN vb_dout0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.960 4.000 81.560 ;
    END
  END vb_dout0[2]
  PIN vb_dout0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 546.080 4.000 546.680 ;
    END
  END vb_dout0[30]
  PIN vb_dout0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 559.680 4.000 560.280 ;
    END
  END vb_dout0[31]
  PIN vb_dout0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 107.480 4.000 108.080 ;
    END
  END vb_dout0[3]
  PIN vb_dout0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 133.320 4.000 133.920 ;
    END
  END vb_dout0[4]
  PIN vb_dout0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 155.760 4.000 156.360 ;
    END
  END vb_dout0[5]
  PIN vb_dout0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 177.520 4.000 178.120 ;
    END
  END vb_dout0[6]
  PIN vb_dout0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 199.280 4.000 199.880 ;
    END
  END vb_dout0[7]
  PIN vb_dout0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 221.040 4.000 221.640 ;
    END
  END vb_dout0[8]
  PIN vb_dout0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 243.480 4.000 244.080 ;
    END
  END vb_dout0[9]
  PIN vb_dout1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.680 4.000 33.280 ;
    END
  END vb_dout1[0]
  PIN vb_dout1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 270.000 4.000 270.600 ;
    END
  END vb_dout1[10]
  PIN vb_dout1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 291.760 4.000 292.360 ;
    END
  END vb_dout1[11]
  PIN vb_dout1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 313.520 4.000 314.120 ;
    END
  END vb_dout1[12]
  PIN vb_dout1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 327.120 4.000 327.720 ;
    END
  END vb_dout1[13]
  PIN vb_dout1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 340.040 4.000 340.640 ;
    END
  END vb_dout1[14]
  PIN vb_dout1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 352.960 4.000 353.560 ;
    END
  END vb_dout1[15]
  PIN vb_dout1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 366.560 4.000 367.160 ;
    END
  END vb_dout1[16]
  PIN vb_dout1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 379.480 4.000 380.080 ;
    END
  END vb_dout1[17]
  PIN vb_dout1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 392.400 4.000 393.000 ;
    END
  END vb_dout1[18]
  PIN vb_dout1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 406.000 4.000 406.600 ;
    END
  END vb_dout1[19]
  PIN vb_dout1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 58.520 4.000 59.120 ;
    END
  END vb_dout1[1]
  PIN vb_dout1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 418.920 4.000 419.520 ;
    END
  END vb_dout1[20]
  PIN vb_dout1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 432.520 4.000 433.120 ;
    END
  END vb_dout1[21]
  PIN vb_dout1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 445.440 4.000 446.040 ;
    END
  END vb_dout1[22]
  PIN vb_dout1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 458.360 4.000 458.960 ;
    END
  END vb_dout1[23]
  PIN vb_dout1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 471.960 4.000 472.560 ;
    END
  END vb_dout1[24]
  PIN vb_dout1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 484.880 4.000 485.480 ;
    END
  END vb_dout1[25]
  PIN vb_dout1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 497.800 4.000 498.400 ;
    END
  END vb_dout1[26]
  PIN vb_dout1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 511.400 4.000 512.000 ;
    END
  END vb_dout1[27]
  PIN vb_dout1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 524.320 4.000 524.920 ;
    END
  END vb_dout1[28]
  PIN vb_dout1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 537.920 4.000 538.520 ;
    END
  END vb_dout1[29]
  PIN vb_dout1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.040 4.000 85.640 ;
    END
  END vb_dout1[2]
  PIN vb_dout1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 550.840 4.000 551.440 ;
    END
  END vb_dout1[30]
  PIN vb_dout1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 563.760 4.000 564.360 ;
    END
  END vb_dout1[31]
  PIN vb_dout1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 111.560 4.000 112.160 ;
    END
  END vb_dout1[3]
  PIN vb_dout1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 138.080 4.000 138.680 ;
    END
  END vb_dout1[4]
  PIN vb_dout1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.840 4.000 160.440 ;
    END
  END vb_dout1[5]
  PIN vb_dout1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 181.600 4.000 182.200 ;
    END
  END vb_dout1[6]
  PIN vb_dout1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.040 4.000 204.640 ;
    END
  END vb_dout1[7]
  PIN vb_dout1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 225.800 4.000 226.400 ;
    END
  END vb_dout1[8]
  PIN vb_dout1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 247.560 4.000 248.160 ;
    END
  END vb_dout1[9]
  PIN vb_web0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.240 4.000 10.840 ;
    END
  END vb_web0
  PIN vb_wmask0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.760 4.000 37.360 ;
    END
  END vb_wmask0[0]
  PIN vb_wmask0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.280 4.000 63.880 ;
    END
  END vb_wmask0[1]
  PIN vb_wmask0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.800 4.000 90.400 ;
    END
  END vb_wmask0[2]
  PIN vb_wmask0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 4.000 116.240 ;
    END
  END vb_wmask0[3]
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1286.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 1286.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 1286.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 1286.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 1286.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 1286.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 1286.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 1286.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.840 10.640 1251.440 1286.800 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 1286.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 1286.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 1286.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 1286.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 1286.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 1286.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 1286.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 1286.800 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 1294.440 1286.645 ;
      LAYER met1 ;
        RECT 2.830 9.900 1294.440 1286.800 ;
      LAYER met2 ;
        RECT 2.860 4.280 1291.120 1297.965 ;
        RECT 2.860 2.195 8.090 4.280 ;
        RECT 8.930 2.195 25.110 4.280 ;
        RECT 25.950 2.195 42.590 4.280 ;
        RECT 43.430 2.195 60.070 4.280 ;
        RECT 60.910 2.195 77.090 4.280 ;
        RECT 77.930 2.195 94.570 4.280 ;
        RECT 95.410 2.195 112.050 4.280 ;
        RECT 112.890 2.195 129.070 4.280 ;
        RECT 129.910 2.195 146.550 4.280 ;
        RECT 147.390 2.195 164.030 4.280 ;
        RECT 164.870 2.195 181.050 4.280 ;
        RECT 181.890 2.195 198.530 4.280 ;
        RECT 199.370 2.195 216.010 4.280 ;
        RECT 216.850 2.195 233.030 4.280 ;
        RECT 233.870 2.195 250.510 4.280 ;
        RECT 251.350 2.195 267.990 4.280 ;
        RECT 268.830 2.195 285.010 4.280 ;
        RECT 285.850 2.195 302.490 4.280 ;
        RECT 303.330 2.195 319.970 4.280 ;
        RECT 320.810 2.195 336.990 4.280 ;
        RECT 337.830 2.195 354.470 4.280 ;
        RECT 355.310 2.195 371.950 4.280 ;
        RECT 372.790 2.195 388.970 4.280 ;
        RECT 389.810 2.195 406.450 4.280 ;
        RECT 407.290 2.195 423.930 4.280 ;
        RECT 424.770 2.195 441.410 4.280 ;
        RECT 442.250 2.195 458.430 4.280 ;
        RECT 459.270 2.195 475.910 4.280 ;
        RECT 476.750 2.195 493.390 4.280 ;
        RECT 494.230 2.195 510.410 4.280 ;
        RECT 511.250 2.195 527.890 4.280 ;
        RECT 528.730 2.195 545.370 4.280 ;
        RECT 546.210 2.195 562.390 4.280 ;
        RECT 563.230 2.195 579.870 4.280 ;
        RECT 580.710 2.195 597.350 4.280 ;
        RECT 598.190 2.195 614.370 4.280 ;
        RECT 615.210 2.195 631.850 4.280 ;
        RECT 632.690 2.195 649.330 4.280 ;
        RECT 650.170 2.195 666.350 4.280 ;
        RECT 667.190 2.195 683.830 4.280 ;
        RECT 684.670 2.195 701.310 4.280 ;
        RECT 702.150 2.195 718.330 4.280 ;
        RECT 719.170 2.195 735.810 4.280 ;
        RECT 736.650 2.195 753.290 4.280 ;
        RECT 754.130 2.195 770.310 4.280 ;
        RECT 771.150 2.195 787.790 4.280 ;
        RECT 788.630 2.195 805.270 4.280 ;
        RECT 806.110 2.195 822.290 4.280 ;
        RECT 823.130 2.195 839.770 4.280 ;
        RECT 840.610 2.195 857.250 4.280 ;
        RECT 858.090 2.195 874.730 4.280 ;
        RECT 875.570 2.195 891.750 4.280 ;
        RECT 892.590 2.195 909.230 4.280 ;
        RECT 910.070 2.195 926.710 4.280 ;
        RECT 927.550 2.195 943.730 4.280 ;
        RECT 944.570 2.195 961.210 4.280 ;
        RECT 962.050 2.195 978.690 4.280 ;
        RECT 979.530 2.195 995.710 4.280 ;
        RECT 996.550 2.195 1013.190 4.280 ;
        RECT 1014.030 2.195 1030.670 4.280 ;
        RECT 1031.510 2.195 1047.690 4.280 ;
        RECT 1048.530 2.195 1065.170 4.280 ;
        RECT 1066.010 2.195 1082.650 4.280 ;
        RECT 1083.490 2.195 1099.670 4.280 ;
        RECT 1100.510 2.195 1117.150 4.280 ;
        RECT 1117.990 2.195 1134.630 4.280 ;
        RECT 1135.470 2.195 1151.650 4.280 ;
        RECT 1152.490 2.195 1169.130 4.280 ;
        RECT 1169.970 2.195 1186.610 4.280 ;
        RECT 1187.450 2.195 1203.630 4.280 ;
        RECT 1204.470 2.195 1221.110 4.280 ;
        RECT 1221.950 2.195 1238.590 4.280 ;
        RECT 1239.430 2.195 1255.610 4.280 ;
        RECT 1256.450 2.195 1273.090 4.280 ;
        RECT 1273.930 2.195 1290.570 4.280 ;
      LAYER met3 ;
        RECT 4.400 1297.080 1251.440 1297.945 ;
        RECT 3.030 1294.400 1251.440 1297.080 ;
        RECT 4.400 1293.000 1251.440 1294.400 ;
        RECT 3.030 1289.640 1251.440 1293.000 ;
        RECT 4.400 1288.240 1251.440 1289.640 ;
        RECT 3.030 1285.560 1251.440 1288.240 ;
        RECT 4.400 1284.160 1251.440 1285.560 ;
        RECT 3.030 1280.800 1251.440 1284.160 ;
        RECT 4.400 1279.400 1251.440 1280.800 ;
        RECT 3.030 1276.720 1251.440 1279.400 ;
        RECT 4.400 1275.320 1251.440 1276.720 ;
        RECT 3.030 1271.960 1251.440 1275.320 ;
        RECT 4.400 1270.560 1251.440 1271.960 ;
        RECT 3.030 1267.880 1251.440 1270.560 ;
        RECT 4.400 1266.480 1251.440 1267.880 ;
        RECT 3.030 1263.120 1251.440 1266.480 ;
        RECT 4.400 1261.720 1251.440 1263.120 ;
        RECT 3.030 1259.040 1251.440 1261.720 ;
        RECT 4.400 1257.640 1251.440 1259.040 ;
        RECT 3.030 1254.280 1251.440 1257.640 ;
        RECT 4.400 1252.880 1251.440 1254.280 ;
        RECT 3.030 1250.200 1251.440 1252.880 ;
        RECT 4.400 1248.800 1251.440 1250.200 ;
        RECT 3.030 1246.120 1251.440 1248.800 ;
        RECT 4.400 1244.720 1251.440 1246.120 ;
        RECT 3.030 1241.360 1251.440 1244.720 ;
        RECT 4.400 1239.960 1251.440 1241.360 ;
        RECT 3.030 1237.280 1251.440 1239.960 ;
        RECT 4.400 1235.880 1251.440 1237.280 ;
        RECT 3.030 1232.520 1251.440 1235.880 ;
        RECT 4.400 1231.120 1251.440 1232.520 ;
        RECT 3.030 1228.440 1251.440 1231.120 ;
        RECT 4.400 1227.040 1251.440 1228.440 ;
        RECT 3.030 1223.680 1251.440 1227.040 ;
        RECT 4.400 1222.280 1251.440 1223.680 ;
        RECT 3.030 1219.600 1251.440 1222.280 ;
        RECT 4.400 1218.200 1251.440 1219.600 ;
        RECT 3.030 1214.840 1251.440 1218.200 ;
        RECT 4.400 1213.440 1251.440 1214.840 ;
        RECT 3.030 1210.760 1251.440 1213.440 ;
        RECT 4.400 1209.360 1251.440 1210.760 ;
        RECT 3.030 1206.000 1251.440 1209.360 ;
        RECT 4.400 1204.600 1251.440 1206.000 ;
        RECT 3.030 1201.920 1251.440 1204.600 ;
        RECT 4.400 1200.520 1251.440 1201.920 ;
        RECT 3.030 1197.160 1251.440 1200.520 ;
        RECT 4.400 1195.760 1251.440 1197.160 ;
        RECT 3.030 1193.080 1251.440 1195.760 ;
        RECT 4.400 1191.680 1251.440 1193.080 ;
        RECT 3.030 1189.000 1251.440 1191.680 ;
        RECT 4.400 1187.600 1251.440 1189.000 ;
        RECT 3.030 1184.240 1251.440 1187.600 ;
        RECT 4.400 1182.840 1251.440 1184.240 ;
        RECT 3.030 1180.160 1251.440 1182.840 ;
        RECT 4.400 1178.760 1251.440 1180.160 ;
        RECT 3.030 1175.400 1251.440 1178.760 ;
        RECT 4.400 1174.000 1251.440 1175.400 ;
        RECT 3.030 1171.320 1251.440 1174.000 ;
        RECT 4.400 1169.920 1251.440 1171.320 ;
        RECT 3.030 1166.560 1251.440 1169.920 ;
        RECT 4.400 1165.160 1251.440 1166.560 ;
        RECT 3.030 1162.480 1251.440 1165.160 ;
        RECT 4.400 1161.080 1251.440 1162.480 ;
        RECT 3.030 1157.720 1251.440 1161.080 ;
        RECT 4.400 1156.320 1251.440 1157.720 ;
        RECT 3.030 1153.640 1251.440 1156.320 ;
        RECT 4.400 1152.240 1251.440 1153.640 ;
        RECT 3.030 1148.880 1251.440 1152.240 ;
        RECT 4.400 1147.480 1251.440 1148.880 ;
        RECT 3.030 1144.800 1251.440 1147.480 ;
        RECT 4.400 1143.400 1251.440 1144.800 ;
        RECT 3.030 1140.720 1251.440 1143.400 ;
        RECT 4.400 1139.320 1251.440 1140.720 ;
        RECT 3.030 1135.960 1251.440 1139.320 ;
        RECT 4.400 1134.560 1251.440 1135.960 ;
        RECT 3.030 1131.880 1251.440 1134.560 ;
        RECT 4.400 1130.480 1251.440 1131.880 ;
        RECT 3.030 1127.120 1251.440 1130.480 ;
        RECT 4.400 1125.720 1251.440 1127.120 ;
        RECT 3.030 1123.040 1251.440 1125.720 ;
        RECT 4.400 1121.640 1251.440 1123.040 ;
        RECT 3.030 1118.280 1251.440 1121.640 ;
        RECT 4.400 1116.880 1251.440 1118.280 ;
        RECT 3.030 1114.200 1251.440 1116.880 ;
        RECT 4.400 1112.800 1251.440 1114.200 ;
        RECT 3.030 1109.440 1251.440 1112.800 ;
        RECT 4.400 1108.040 1251.440 1109.440 ;
        RECT 3.030 1105.360 1251.440 1108.040 ;
        RECT 4.400 1103.960 1251.440 1105.360 ;
        RECT 3.030 1100.600 1251.440 1103.960 ;
        RECT 4.400 1099.200 1251.440 1100.600 ;
        RECT 3.030 1096.520 1251.440 1099.200 ;
        RECT 4.400 1095.120 1251.440 1096.520 ;
        RECT 3.030 1091.760 1251.440 1095.120 ;
        RECT 4.400 1090.360 1251.440 1091.760 ;
        RECT 3.030 1087.680 1251.440 1090.360 ;
        RECT 4.400 1086.280 1251.440 1087.680 ;
        RECT 3.030 1083.600 1251.440 1086.280 ;
        RECT 4.400 1082.200 1251.440 1083.600 ;
        RECT 3.030 1078.840 1251.440 1082.200 ;
        RECT 4.400 1077.440 1251.440 1078.840 ;
        RECT 3.030 1074.760 1251.440 1077.440 ;
        RECT 4.400 1073.360 1251.440 1074.760 ;
        RECT 3.030 1070.000 1251.440 1073.360 ;
        RECT 4.400 1068.600 1251.440 1070.000 ;
        RECT 3.030 1065.920 1251.440 1068.600 ;
        RECT 4.400 1064.520 1251.440 1065.920 ;
        RECT 3.030 1061.160 1251.440 1064.520 ;
        RECT 4.400 1059.760 1251.440 1061.160 ;
        RECT 3.030 1057.080 1251.440 1059.760 ;
        RECT 4.400 1055.680 1251.440 1057.080 ;
        RECT 3.030 1052.320 1251.440 1055.680 ;
        RECT 4.400 1050.920 1251.440 1052.320 ;
        RECT 3.030 1048.240 1251.440 1050.920 ;
        RECT 4.400 1046.840 1251.440 1048.240 ;
        RECT 3.030 1043.480 1251.440 1046.840 ;
        RECT 4.400 1042.080 1251.440 1043.480 ;
        RECT 3.030 1039.400 1251.440 1042.080 ;
        RECT 4.400 1038.000 1251.440 1039.400 ;
        RECT 3.030 1034.640 1251.440 1038.000 ;
        RECT 4.400 1033.240 1251.440 1034.640 ;
        RECT 3.030 1030.560 1251.440 1033.240 ;
        RECT 4.400 1029.160 1251.440 1030.560 ;
        RECT 3.030 1026.480 1251.440 1029.160 ;
        RECT 4.400 1025.080 1251.440 1026.480 ;
        RECT 3.030 1021.720 1251.440 1025.080 ;
        RECT 4.400 1020.320 1251.440 1021.720 ;
        RECT 3.030 1017.640 1251.440 1020.320 ;
        RECT 4.400 1016.240 1251.440 1017.640 ;
        RECT 3.030 1012.880 1251.440 1016.240 ;
        RECT 4.400 1011.480 1251.440 1012.880 ;
        RECT 3.030 1008.800 1251.440 1011.480 ;
        RECT 4.400 1007.400 1251.440 1008.800 ;
        RECT 3.030 1004.040 1251.440 1007.400 ;
        RECT 4.400 1002.640 1251.440 1004.040 ;
        RECT 3.030 999.960 1251.440 1002.640 ;
        RECT 4.400 998.560 1251.440 999.960 ;
        RECT 3.030 995.200 1251.440 998.560 ;
        RECT 4.400 993.800 1251.440 995.200 ;
        RECT 3.030 991.120 1251.440 993.800 ;
        RECT 4.400 989.720 1251.440 991.120 ;
        RECT 3.030 986.360 1251.440 989.720 ;
        RECT 4.400 984.960 1251.440 986.360 ;
        RECT 3.030 982.280 1251.440 984.960 ;
        RECT 4.400 980.880 1251.440 982.280 ;
        RECT 3.030 978.200 1251.440 980.880 ;
        RECT 4.400 976.800 1251.440 978.200 ;
        RECT 3.030 973.440 1251.440 976.800 ;
        RECT 4.400 972.040 1251.440 973.440 ;
        RECT 3.030 969.360 1251.440 972.040 ;
        RECT 4.400 967.960 1251.440 969.360 ;
        RECT 3.030 964.600 1251.440 967.960 ;
        RECT 4.400 963.200 1251.440 964.600 ;
        RECT 3.030 960.520 1251.440 963.200 ;
        RECT 4.400 959.120 1251.440 960.520 ;
        RECT 3.030 955.760 1251.440 959.120 ;
        RECT 4.400 954.360 1251.440 955.760 ;
        RECT 3.030 951.680 1251.440 954.360 ;
        RECT 4.400 950.280 1251.440 951.680 ;
        RECT 3.030 946.920 1251.440 950.280 ;
        RECT 4.400 945.520 1251.440 946.920 ;
        RECT 3.030 942.840 1251.440 945.520 ;
        RECT 4.400 941.440 1251.440 942.840 ;
        RECT 3.030 938.080 1251.440 941.440 ;
        RECT 4.400 936.680 1251.440 938.080 ;
        RECT 3.030 934.000 1251.440 936.680 ;
        RECT 4.400 932.600 1251.440 934.000 ;
        RECT 3.030 929.240 1251.440 932.600 ;
        RECT 4.400 927.840 1251.440 929.240 ;
        RECT 3.030 925.160 1251.440 927.840 ;
        RECT 4.400 923.760 1251.440 925.160 ;
        RECT 3.030 921.080 1251.440 923.760 ;
        RECT 4.400 919.680 1251.440 921.080 ;
        RECT 3.030 916.320 1251.440 919.680 ;
        RECT 4.400 914.920 1251.440 916.320 ;
        RECT 3.030 912.240 1251.440 914.920 ;
        RECT 4.400 910.840 1251.440 912.240 ;
        RECT 3.030 907.480 1251.440 910.840 ;
        RECT 4.400 906.080 1251.440 907.480 ;
        RECT 3.030 903.400 1251.440 906.080 ;
        RECT 4.400 902.000 1251.440 903.400 ;
        RECT 3.030 898.640 1251.440 902.000 ;
        RECT 4.400 897.240 1251.440 898.640 ;
        RECT 3.030 894.560 1251.440 897.240 ;
        RECT 4.400 893.160 1251.440 894.560 ;
        RECT 3.030 889.800 1251.440 893.160 ;
        RECT 4.400 888.400 1251.440 889.800 ;
        RECT 3.030 885.720 1251.440 888.400 ;
        RECT 4.400 884.320 1251.440 885.720 ;
        RECT 3.030 880.960 1251.440 884.320 ;
        RECT 4.400 879.560 1251.440 880.960 ;
        RECT 3.030 876.880 1251.440 879.560 ;
        RECT 4.400 875.480 1251.440 876.880 ;
        RECT 3.030 872.120 1251.440 875.480 ;
        RECT 4.400 870.720 1251.440 872.120 ;
        RECT 3.030 868.040 1251.440 870.720 ;
        RECT 4.400 866.640 1251.440 868.040 ;
        RECT 3.030 863.960 1251.440 866.640 ;
        RECT 4.400 862.560 1251.440 863.960 ;
        RECT 3.030 859.200 1251.440 862.560 ;
        RECT 4.400 857.800 1251.440 859.200 ;
        RECT 3.030 855.120 1251.440 857.800 ;
        RECT 4.400 853.720 1251.440 855.120 ;
        RECT 3.030 850.360 1251.440 853.720 ;
        RECT 4.400 848.960 1251.440 850.360 ;
        RECT 3.030 846.280 1251.440 848.960 ;
        RECT 4.400 844.880 1251.440 846.280 ;
        RECT 3.030 841.520 1251.440 844.880 ;
        RECT 4.400 840.120 1251.440 841.520 ;
        RECT 3.030 837.440 1251.440 840.120 ;
        RECT 4.400 836.040 1251.440 837.440 ;
        RECT 3.030 832.680 1251.440 836.040 ;
        RECT 4.400 831.280 1251.440 832.680 ;
        RECT 3.030 828.600 1251.440 831.280 ;
        RECT 4.400 827.200 1251.440 828.600 ;
        RECT 3.030 823.840 1251.440 827.200 ;
        RECT 4.400 822.440 1251.440 823.840 ;
        RECT 3.030 819.760 1251.440 822.440 ;
        RECT 4.400 818.360 1251.440 819.760 ;
        RECT 3.030 815.680 1251.440 818.360 ;
        RECT 4.400 814.280 1251.440 815.680 ;
        RECT 3.030 810.920 1251.440 814.280 ;
        RECT 4.400 809.520 1251.440 810.920 ;
        RECT 3.030 806.840 1251.440 809.520 ;
        RECT 4.400 805.440 1251.440 806.840 ;
        RECT 3.030 802.080 1251.440 805.440 ;
        RECT 4.400 800.680 1251.440 802.080 ;
        RECT 3.030 798.000 1251.440 800.680 ;
        RECT 4.400 796.600 1251.440 798.000 ;
        RECT 3.030 793.240 1251.440 796.600 ;
        RECT 4.400 791.840 1251.440 793.240 ;
        RECT 3.030 789.160 1251.440 791.840 ;
        RECT 4.400 787.760 1251.440 789.160 ;
        RECT 3.030 784.400 1251.440 787.760 ;
        RECT 4.400 783.000 1251.440 784.400 ;
        RECT 3.030 780.320 1251.440 783.000 ;
        RECT 4.400 778.920 1251.440 780.320 ;
        RECT 3.030 775.560 1251.440 778.920 ;
        RECT 4.400 774.160 1251.440 775.560 ;
        RECT 3.030 771.480 1251.440 774.160 ;
        RECT 4.400 770.080 1251.440 771.480 ;
        RECT 3.030 766.720 1251.440 770.080 ;
        RECT 4.400 765.320 1251.440 766.720 ;
        RECT 3.030 762.640 1251.440 765.320 ;
        RECT 4.400 761.240 1251.440 762.640 ;
        RECT 3.030 758.560 1251.440 761.240 ;
        RECT 4.400 757.160 1251.440 758.560 ;
        RECT 3.030 753.800 1251.440 757.160 ;
        RECT 4.400 752.400 1251.440 753.800 ;
        RECT 3.030 749.720 1251.440 752.400 ;
        RECT 4.400 748.320 1251.440 749.720 ;
        RECT 3.030 744.960 1251.440 748.320 ;
        RECT 4.400 743.560 1251.440 744.960 ;
        RECT 3.030 740.880 1251.440 743.560 ;
        RECT 4.400 739.480 1251.440 740.880 ;
        RECT 3.030 736.120 1251.440 739.480 ;
        RECT 4.400 734.720 1251.440 736.120 ;
        RECT 3.030 732.040 1251.440 734.720 ;
        RECT 4.400 730.640 1251.440 732.040 ;
        RECT 3.030 727.280 1251.440 730.640 ;
        RECT 4.400 725.880 1251.440 727.280 ;
        RECT 3.030 723.200 1251.440 725.880 ;
        RECT 4.400 721.800 1251.440 723.200 ;
        RECT 3.030 718.440 1251.440 721.800 ;
        RECT 4.400 717.040 1251.440 718.440 ;
        RECT 3.030 714.360 1251.440 717.040 ;
        RECT 4.400 712.960 1251.440 714.360 ;
        RECT 3.030 709.600 1251.440 712.960 ;
        RECT 4.400 708.200 1251.440 709.600 ;
        RECT 3.030 705.520 1251.440 708.200 ;
        RECT 4.400 704.120 1251.440 705.520 ;
        RECT 3.030 701.440 1251.440 704.120 ;
        RECT 4.400 700.040 1251.440 701.440 ;
        RECT 3.030 696.680 1251.440 700.040 ;
        RECT 4.400 695.280 1251.440 696.680 ;
        RECT 3.030 692.600 1251.440 695.280 ;
        RECT 4.400 691.200 1251.440 692.600 ;
        RECT 3.030 687.840 1251.440 691.200 ;
        RECT 4.400 686.440 1251.440 687.840 ;
        RECT 3.030 683.760 1251.440 686.440 ;
        RECT 4.400 682.360 1251.440 683.760 ;
        RECT 3.030 679.000 1251.440 682.360 ;
        RECT 4.400 677.600 1251.440 679.000 ;
        RECT 3.030 674.920 1251.440 677.600 ;
        RECT 4.400 673.520 1251.440 674.920 ;
        RECT 3.030 670.160 1251.440 673.520 ;
        RECT 4.400 668.760 1251.440 670.160 ;
        RECT 3.030 666.080 1251.440 668.760 ;
        RECT 4.400 664.680 1251.440 666.080 ;
        RECT 3.030 661.320 1251.440 664.680 ;
        RECT 4.400 659.920 1251.440 661.320 ;
        RECT 3.030 657.240 1251.440 659.920 ;
        RECT 4.400 655.840 1251.440 657.240 ;
        RECT 3.030 653.160 1251.440 655.840 ;
        RECT 4.400 651.760 1251.440 653.160 ;
        RECT 3.030 648.400 1251.440 651.760 ;
        RECT 4.400 647.000 1251.440 648.400 ;
        RECT 3.030 644.320 1251.440 647.000 ;
        RECT 4.400 642.920 1251.440 644.320 ;
        RECT 3.030 639.560 1251.440 642.920 ;
        RECT 4.400 638.160 1251.440 639.560 ;
        RECT 3.030 635.480 1251.440 638.160 ;
        RECT 4.400 634.080 1251.440 635.480 ;
        RECT 3.030 630.720 1251.440 634.080 ;
        RECT 4.400 629.320 1251.440 630.720 ;
        RECT 3.030 626.640 1251.440 629.320 ;
        RECT 4.400 625.240 1251.440 626.640 ;
        RECT 3.030 621.880 1251.440 625.240 ;
        RECT 4.400 620.480 1251.440 621.880 ;
        RECT 3.030 617.800 1251.440 620.480 ;
        RECT 4.400 616.400 1251.440 617.800 ;
        RECT 3.030 613.040 1251.440 616.400 ;
        RECT 4.400 611.640 1251.440 613.040 ;
        RECT 3.030 608.960 1251.440 611.640 ;
        RECT 4.400 607.560 1251.440 608.960 ;
        RECT 3.030 604.200 1251.440 607.560 ;
        RECT 4.400 602.800 1251.440 604.200 ;
        RECT 3.030 600.120 1251.440 602.800 ;
        RECT 4.400 598.720 1251.440 600.120 ;
        RECT 3.030 596.040 1251.440 598.720 ;
        RECT 4.400 594.640 1251.440 596.040 ;
        RECT 3.030 591.280 1251.440 594.640 ;
        RECT 4.400 589.880 1251.440 591.280 ;
        RECT 3.030 587.200 1251.440 589.880 ;
        RECT 4.400 585.800 1251.440 587.200 ;
        RECT 3.030 582.440 1251.440 585.800 ;
        RECT 4.400 581.040 1251.440 582.440 ;
        RECT 3.030 578.360 1251.440 581.040 ;
        RECT 4.400 576.960 1251.440 578.360 ;
        RECT 3.030 573.600 1251.440 576.960 ;
        RECT 4.400 572.200 1251.440 573.600 ;
        RECT 3.030 569.520 1251.440 572.200 ;
        RECT 4.400 568.120 1251.440 569.520 ;
        RECT 3.030 564.760 1251.440 568.120 ;
        RECT 4.400 563.360 1251.440 564.760 ;
        RECT 3.030 560.680 1251.440 563.360 ;
        RECT 4.400 559.280 1251.440 560.680 ;
        RECT 3.030 555.920 1251.440 559.280 ;
        RECT 4.400 554.520 1251.440 555.920 ;
        RECT 3.030 551.840 1251.440 554.520 ;
        RECT 4.400 550.440 1251.440 551.840 ;
        RECT 3.030 547.080 1251.440 550.440 ;
        RECT 4.400 545.680 1251.440 547.080 ;
        RECT 3.030 543.000 1251.440 545.680 ;
        RECT 4.400 541.600 1251.440 543.000 ;
        RECT 3.030 538.920 1251.440 541.600 ;
        RECT 4.400 537.520 1251.440 538.920 ;
        RECT 3.030 534.160 1251.440 537.520 ;
        RECT 4.400 532.760 1251.440 534.160 ;
        RECT 3.030 530.080 1251.440 532.760 ;
        RECT 4.400 528.680 1251.440 530.080 ;
        RECT 3.030 525.320 1251.440 528.680 ;
        RECT 4.400 523.920 1251.440 525.320 ;
        RECT 3.030 521.240 1251.440 523.920 ;
        RECT 4.400 519.840 1251.440 521.240 ;
        RECT 3.030 516.480 1251.440 519.840 ;
        RECT 4.400 515.080 1251.440 516.480 ;
        RECT 3.030 512.400 1251.440 515.080 ;
        RECT 4.400 511.000 1251.440 512.400 ;
        RECT 3.030 507.640 1251.440 511.000 ;
        RECT 4.400 506.240 1251.440 507.640 ;
        RECT 3.030 503.560 1251.440 506.240 ;
        RECT 4.400 502.160 1251.440 503.560 ;
        RECT 3.030 498.800 1251.440 502.160 ;
        RECT 4.400 497.400 1251.440 498.800 ;
        RECT 3.030 494.720 1251.440 497.400 ;
        RECT 4.400 493.320 1251.440 494.720 ;
        RECT 3.030 490.640 1251.440 493.320 ;
        RECT 4.400 489.240 1251.440 490.640 ;
        RECT 3.030 485.880 1251.440 489.240 ;
        RECT 4.400 484.480 1251.440 485.880 ;
        RECT 3.030 481.800 1251.440 484.480 ;
        RECT 4.400 480.400 1251.440 481.800 ;
        RECT 3.030 477.040 1251.440 480.400 ;
        RECT 4.400 475.640 1251.440 477.040 ;
        RECT 3.030 472.960 1251.440 475.640 ;
        RECT 4.400 471.560 1251.440 472.960 ;
        RECT 3.030 468.200 1251.440 471.560 ;
        RECT 4.400 466.800 1251.440 468.200 ;
        RECT 3.030 464.120 1251.440 466.800 ;
        RECT 4.400 462.720 1251.440 464.120 ;
        RECT 3.030 459.360 1251.440 462.720 ;
        RECT 4.400 457.960 1251.440 459.360 ;
        RECT 3.030 455.280 1251.440 457.960 ;
        RECT 4.400 453.880 1251.440 455.280 ;
        RECT 3.030 450.520 1251.440 453.880 ;
        RECT 4.400 449.120 1251.440 450.520 ;
        RECT 3.030 446.440 1251.440 449.120 ;
        RECT 4.400 445.040 1251.440 446.440 ;
        RECT 3.030 441.680 1251.440 445.040 ;
        RECT 4.400 440.280 1251.440 441.680 ;
        RECT 3.030 437.600 1251.440 440.280 ;
        RECT 4.400 436.200 1251.440 437.600 ;
        RECT 3.030 433.520 1251.440 436.200 ;
        RECT 4.400 432.120 1251.440 433.520 ;
        RECT 3.030 428.760 1251.440 432.120 ;
        RECT 4.400 427.360 1251.440 428.760 ;
        RECT 3.030 424.680 1251.440 427.360 ;
        RECT 4.400 423.280 1251.440 424.680 ;
        RECT 3.030 419.920 1251.440 423.280 ;
        RECT 4.400 418.520 1251.440 419.920 ;
        RECT 3.030 415.840 1251.440 418.520 ;
        RECT 4.400 414.440 1251.440 415.840 ;
        RECT 3.030 411.080 1251.440 414.440 ;
        RECT 4.400 409.680 1251.440 411.080 ;
        RECT 3.030 407.000 1251.440 409.680 ;
        RECT 4.400 405.600 1251.440 407.000 ;
        RECT 3.030 402.240 1251.440 405.600 ;
        RECT 4.400 400.840 1251.440 402.240 ;
        RECT 3.030 398.160 1251.440 400.840 ;
        RECT 4.400 396.760 1251.440 398.160 ;
        RECT 3.030 393.400 1251.440 396.760 ;
        RECT 4.400 392.000 1251.440 393.400 ;
        RECT 3.030 389.320 1251.440 392.000 ;
        RECT 4.400 387.920 1251.440 389.320 ;
        RECT 3.030 384.560 1251.440 387.920 ;
        RECT 4.400 383.160 1251.440 384.560 ;
        RECT 3.030 380.480 1251.440 383.160 ;
        RECT 4.400 379.080 1251.440 380.480 ;
        RECT 3.030 376.400 1251.440 379.080 ;
        RECT 4.400 375.000 1251.440 376.400 ;
        RECT 3.030 371.640 1251.440 375.000 ;
        RECT 4.400 370.240 1251.440 371.640 ;
        RECT 3.030 367.560 1251.440 370.240 ;
        RECT 4.400 366.160 1251.440 367.560 ;
        RECT 3.030 362.800 1251.440 366.160 ;
        RECT 4.400 361.400 1251.440 362.800 ;
        RECT 3.030 358.720 1251.440 361.400 ;
        RECT 4.400 357.320 1251.440 358.720 ;
        RECT 3.030 353.960 1251.440 357.320 ;
        RECT 4.400 352.560 1251.440 353.960 ;
        RECT 3.030 349.880 1251.440 352.560 ;
        RECT 4.400 348.480 1251.440 349.880 ;
        RECT 3.030 345.120 1251.440 348.480 ;
        RECT 4.400 343.720 1251.440 345.120 ;
        RECT 3.030 341.040 1251.440 343.720 ;
        RECT 4.400 339.640 1251.440 341.040 ;
        RECT 3.030 336.280 1251.440 339.640 ;
        RECT 4.400 334.880 1251.440 336.280 ;
        RECT 3.030 332.200 1251.440 334.880 ;
        RECT 4.400 330.800 1251.440 332.200 ;
        RECT 3.030 328.120 1251.440 330.800 ;
        RECT 4.400 326.720 1251.440 328.120 ;
        RECT 3.030 323.360 1251.440 326.720 ;
        RECT 4.400 321.960 1251.440 323.360 ;
        RECT 3.030 319.280 1251.440 321.960 ;
        RECT 4.400 317.880 1251.440 319.280 ;
        RECT 3.030 314.520 1251.440 317.880 ;
        RECT 4.400 313.120 1251.440 314.520 ;
        RECT 3.030 310.440 1251.440 313.120 ;
        RECT 4.400 309.040 1251.440 310.440 ;
        RECT 3.030 305.680 1251.440 309.040 ;
        RECT 4.400 304.280 1251.440 305.680 ;
        RECT 3.030 301.600 1251.440 304.280 ;
        RECT 4.400 300.200 1251.440 301.600 ;
        RECT 3.030 296.840 1251.440 300.200 ;
        RECT 4.400 295.440 1251.440 296.840 ;
        RECT 3.030 292.760 1251.440 295.440 ;
        RECT 4.400 291.360 1251.440 292.760 ;
        RECT 3.030 288.000 1251.440 291.360 ;
        RECT 4.400 286.600 1251.440 288.000 ;
        RECT 3.030 283.920 1251.440 286.600 ;
        RECT 4.400 282.520 1251.440 283.920 ;
        RECT 3.030 279.160 1251.440 282.520 ;
        RECT 4.400 277.760 1251.440 279.160 ;
        RECT 3.030 275.080 1251.440 277.760 ;
        RECT 4.400 273.680 1251.440 275.080 ;
        RECT 3.030 271.000 1251.440 273.680 ;
        RECT 4.400 269.600 1251.440 271.000 ;
        RECT 3.030 266.240 1251.440 269.600 ;
        RECT 4.400 264.840 1251.440 266.240 ;
        RECT 3.030 262.160 1251.440 264.840 ;
        RECT 4.400 260.760 1251.440 262.160 ;
        RECT 3.030 257.400 1251.440 260.760 ;
        RECT 4.400 256.000 1251.440 257.400 ;
        RECT 3.030 253.320 1251.440 256.000 ;
        RECT 4.400 251.920 1251.440 253.320 ;
        RECT 3.030 248.560 1251.440 251.920 ;
        RECT 4.400 247.160 1251.440 248.560 ;
        RECT 3.030 244.480 1251.440 247.160 ;
        RECT 4.400 243.080 1251.440 244.480 ;
        RECT 3.030 239.720 1251.440 243.080 ;
        RECT 4.400 238.320 1251.440 239.720 ;
        RECT 3.030 235.640 1251.440 238.320 ;
        RECT 4.400 234.240 1251.440 235.640 ;
        RECT 3.030 230.880 1251.440 234.240 ;
        RECT 4.400 229.480 1251.440 230.880 ;
        RECT 3.030 226.800 1251.440 229.480 ;
        RECT 4.400 225.400 1251.440 226.800 ;
        RECT 3.030 222.040 1251.440 225.400 ;
        RECT 4.400 220.640 1251.440 222.040 ;
        RECT 3.030 217.960 1251.440 220.640 ;
        RECT 4.400 216.560 1251.440 217.960 ;
        RECT 3.030 213.880 1251.440 216.560 ;
        RECT 4.400 212.480 1251.440 213.880 ;
        RECT 3.030 209.120 1251.440 212.480 ;
        RECT 4.400 207.720 1251.440 209.120 ;
        RECT 3.030 205.040 1251.440 207.720 ;
        RECT 4.400 203.640 1251.440 205.040 ;
        RECT 3.030 200.280 1251.440 203.640 ;
        RECT 4.400 198.880 1251.440 200.280 ;
        RECT 3.030 196.200 1251.440 198.880 ;
        RECT 4.400 194.800 1251.440 196.200 ;
        RECT 3.030 191.440 1251.440 194.800 ;
        RECT 4.400 190.040 1251.440 191.440 ;
        RECT 3.030 187.360 1251.440 190.040 ;
        RECT 4.400 185.960 1251.440 187.360 ;
        RECT 3.030 182.600 1251.440 185.960 ;
        RECT 4.400 181.200 1251.440 182.600 ;
        RECT 3.030 178.520 1251.440 181.200 ;
        RECT 4.400 177.120 1251.440 178.520 ;
        RECT 3.030 173.760 1251.440 177.120 ;
        RECT 4.400 172.360 1251.440 173.760 ;
        RECT 3.030 169.680 1251.440 172.360 ;
        RECT 4.400 168.280 1251.440 169.680 ;
        RECT 3.030 165.600 1251.440 168.280 ;
        RECT 4.400 164.200 1251.440 165.600 ;
        RECT 3.030 160.840 1251.440 164.200 ;
        RECT 4.400 159.440 1251.440 160.840 ;
        RECT 3.030 156.760 1251.440 159.440 ;
        RECT 4.400 155.360 1251.440 156.760 ;
        RECT 3.030 152.000 1251.440 155.360 ;
        RECT 4.400 150.600 1251.440 152.000 ;
        RECT 3.030 147.920 1251.440 150.600 ;
        RECT 4.400 146.520 1251.440 147.920 ;
        RECT 3.030 143.160 1251.440 146.520 ;
        RECT 4.400 141.760 1251.440 143.160 ;
        RECT 3.030 139.080 1251.440 141.760 ;
        RECT 4.400 137.680 1251.440 139.080 ;
        RECT 3.030 134.320 1251.440 137.680 ;
        RECT 4.400 132.920 1251.440 134.320 ;
        RECT 3.030 130.240 1251.440 132.920 ;
        RECT 4.400 128.840 1251.440 130.240 ;
        RECT 3.030 125.480 1251.440 128.840 ;
        RECT 4.400 124.080 1251.440 125.480 ;
        RECT 3.030 121.400 1251.440 124.080 ;
        RECT 4.400 120.000 1251.440 121.400 ;
        RECT 3.030 116.640 1251.440 120.000 ;
        RECT 4.400 115.240 1251.440 116.640 ;
        RECT 3.030 112.560 1251.440 115.240 ;
        RECT 4.400 111.160 1251.440 112.560 ;
        RECT 3.030 108.480 1251.440 111.160 ;
        RECT 4.400 107.080 1251.440 108.480 ;
        RECT 3.030 103.720 1251.440 107.080 ;
        RECT 4.400 102.320 1251.440 103.720 ;
        RECT 3.030 99.640 1251.440 102.320 ;
        RECT 4.400 98.240 1251.440 99.640 ;
        RECT 3.030 94.880 1251.440 98.240 ;
        RECT 4.400 93.480 1251.440 94.880 ;
        RECT 3.030 90.800 1251.440 93.480 ;
        RECT 4.400 89.400 1251.440 90.800 ;
        RECT 3.030 86.040 1251.440 89.400 ;
        RECT 4.400 84.640 1251.440 86.040 ;
        RECT 3.030 81.960 1251.440 84.640 ;
        RECT 4.400 80.560 1251.440 81.960 ;
        RECT 3.030 77.200 1251.440 80.560 ;
        RECT 4.400 75.800 1251.440 77.200 ;
        RECT 3.030 73.120 1251.440 75.800 ;
        RECT 4.400 71.720 1251.440 73.120 ;
        RECT 3.030 68.360 1251.440 71.720 ;
        RECT 4.400 66.960 1251.440 68.360 ;
        RECT 3.030 64.280 1251.440 66.960 ;
        RECT 4.400 62.880 1251.440 64.280 ;
        RECT 3.030 59.520 1251.440 62.880 ;
        RECT 4.400 58.120 1251.440 59.520 ;
        RECT 3.030 55.440 1251.440 58.120 ;
        RECT 4.400 54.040 1251.440 55.440 ;
        RECT 3.030 51.360 1251.440 54.040 ;
        RECT 4.400 49.960 1251.440 51.360 ;
        RECT 3.030 46.600 1251.440 49.960 ;
        RECT 4.400 45.200 1251.440 46.600 ;
        RECT 3.030 42.520 1251.440 45.200 ;
        RECT 4.400 41.120 1251.440 42.520 ;
        RECT 3.030 37.760 1251.440 41.120 ;
        RECT 4.400 36.360 1251.440 37.760 ;
        RECT 3.030 33.680 1251.440 36.360 ;
        RECT 4.400 32.280 1251.440 33.680 ;
        RECT 3.030 28.920 1251.440 32.280 ;
        RECT 4.400 27.520 1251.440 28.920 ;
        RECT 3.030 24.840 1251.440 27.520 ;
        RECT 4.400 23.440 1251.440 24.840 ;
        RECT 3.030 20.080 1251.440 23.440 ;
        RECT 4.400 18.680 1251.440 20.080 ;
        RECT 3.030 16.000 1251.440 18.680 ;
        RECT 4.400 14.600 1251.440 16.000 ;
        RECT 3.030 11.240 1251.440 14.600 ;
        RECT 4.400 9.840 1251.440 11.240 ;
        RECT 3.030 7.160 1251.440 9.840 ;
        RECT 4.400 5.760 1251.440 7.160 ;
        RECT 3.030 3.080 1251.440 5.760 ;
        RECT 4.400 2.215 1251.440 3.080 ;
      LAYER met4 ;
        RECT 3.055 11.735 20.640 1273.465 ;
        RECT 23.040 11.735 97.440 1273.465 ;
        RECT 99.840 11.735 174.240 1273.465 ;
        RECT 176.640 11.735 251.040 1273.465 ;
        RECT 253.440 11.735 327.840 1273.465 ;
        RECT 330.240 11.735 404.640 1273.465 ;
        RECT 407.040 11.735 481.440 1273.465 ;
        RECT 483.840 11.735 558.240 1273.465 ;
        RECT 560.640 11.735 635.040 1273.465 ;
        RECT 637.440 11.735 711.840 1273.465 ;
        RECT 714.240 11.735 788.640 1273.465 ;
        RECT 791.040 11.735 865.440 1273.465 ;
        RECT 867.840 11.735 942.240 1273.465 ;
        RECT 944.640 11.735 1011.705 1273.465 ;
  END
END c0_system
END LIBRARY


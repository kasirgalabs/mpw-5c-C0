magic
tech sky130A
magscale 1 2
timestamp 1647616682
<< obsli1 >>
rect 1104 2159 298816 297585
<< obsm1 >>
rect 474 1980 298816 297616
<< metal2 >>
rect 1950 0 2006 800
rect 5906 0 5962 800
rect 9862 0 9918 800
rect 13910 0 13966 800
rect 17866 0 17922 800
rect 21914 0 21970 800
rect 25870 0 25926 800
rect 29918 0 29974 800
rect 33874 0 33930 800
rect 37922 0 37978 800
rect 41878 0 41934 800
rect 45926 0 45982 800
rect 49882 0 49938 800
rect 53930 0 53986 800
rect 57886 0 57942 800
rect 61934 0 61990 800
rect 65890 0 65946 800
rect 69938 0 69994 800
rect 73894 0 73950 800
rect 77942 0 77998 800
rect 81898 0 81954 800
rect 85946 0 86002 800
rect 89902 0 89958 800
rect 93950 0 94006 800
rect 97906 0 97962 800
rect 101954 0 102010 800
rect 105910 0 105966 800
rect 109866 0 109922 800
rect 113914 0 113970 800
rect 117870 0 117926 800
rect 121918 0 121974 800
rect 125874 0 125930 800
rect 129922 0 129978 800
rect 133878 0 133934 800
rect 137926 0 137982 800
rect 141882 0 141938 800
rect 145930 0 145986 800
rect 149886 0 149942 800
rect 153934 0 153990 800
rect 157890 0 157946 800
rect 161938 0 161994 800
rect 165894 0 165950 800
rect 169942 0 169998 800
rect 173898 0 173954 800
rect 177946 0 178002 800
rect 181902 0 181958 800
rect 185950 0 186006 800
rect 189906 0 189962 800
rect 193954 0 194010 800
rect 197910 0 197966 800
rect 201958 0 202014 800
rect 205914 0 205970 800
rect 209870 0 209926 800
rect 213918 0 213974 800
rect 217874 0 217930 800
rect 221922 0 221978 800
rect 225878 0 225934 800
rect 229926 0 229982 800
rect 233882 0 233938 800
rect 237930 0 237986 800
rect 241886 0 241942 800
rect 245934 0 245990 800
rect 249890 0 249946 800
rect 253938 0 253994 800
rect 257894 0 257950 800
rect 261942 0 261998 800
rect 265898 0 265954 800
rect 269946 0 270002 800
rect 273902 0 273958 800
rect 277950 0 278006 800
rect 281906 0 281962 800
rect 285954 0 286010 800
rect 289910 0 289966 800
rect 293958 0 294014 800
rect 297914 0 297970 800
<< obsm2 >>
rect 480 856 297968 299441
rect 480 439 1894 856
rect 2062 439 5850 856
rect 6018 439 9806 856
rect 9974 439 13854 856
rect 14022 439 17810 856
rect 17978 439 21858 856
rect 22026 439 25814 856
rect 25982 439 29862 856
rect 30030 439 33818 856
rect 33986 439 37866 856
rect 38034 439 41822 856
rect 41990 439 45870 856
rect 46038 439 49826 856
rect 49994 439 53874 856
rect 54042 439 57830 856
rect 57998 439 61878 856
rect 62046 439 65834 856
rect 66002 439 69882 856
rect 70050 439 73838 856
rect 74006 439 77886 856
rect 78054 439 81842 856
rect 82010 439 85890 856
rect 86058 439 89846 856
rect 90014 439 93894 856
rect 94062 439 97850 856
rect 98018 439 101898 856
rect 102066 439 105854 856
rect 106022 439 109810 856
rect 109978 439 113858 856
rect 114026 439 117814 856
rect 117982 439 121862 856
rect 122030 439 125818 856
rect 125986 439 129866 856
rect 130034 439 133822 856
rect 133990 439 137870 856
rect 138038 439 141826 856
rect 141994 439 145874 856
rect 146042 439 149830 856
rect 149998 439 153878 856
rect 154046 439 157834 856
rect 158002 439 161882 856
rect 162050 439 165838 856
rect 166006 439 169886 856
rect 170054 439 173842 856
rect 174010 439 177890 856
rect 178058 439 181846 856
rect 182014 439 185894 856
rect 186062 439 189850 856
rect 190018 439 193898 856
rect 194066 439 197854 856
rect 198022 439 201902 856
rect 202070 439 205858 856
rect 206026 439 209814 856
rect 209982 439 213862 856
rect 214030 439 217818 856
rect 217986 439 221866 856
rect 222034 439 225822 856
rect 225990 439 229870 856
rect 230038 439 233826 856
rect 233994 439 237874 856
rect 238042 439 241830 856
rect 241998 439 245878 856
rect 246046 439 249834 856
rect 250002 439 253882 856
rect 254050 439 257838 856
rect 258006 439 261886 856
rect 262054 439 265842 856
rect 266010 439 269890 856
rect 270058 439 273846 856
rect 274014 439 277894 856
rect 278062 439 281850 856
rect 282018 439 285898 856
rect 286066 439 289854 856
rect 290022 439 293902 856
rect 294070 439 297858 856
<< metal3 >>
rect 0 299344 800 299464
rect 0 298392 800 298512
rect 0 297304 800 297424
rect 0 296352 800 296472
rect 0 295264 800 295384
rect 0 294312 800 294432
rect 0 293224 800 293344
rect 0 292272 800 292392
rect 0 291184 800 291304
rect 0 290232 800 290352
rect 0 289280 800 289400
rect 0 288192 800 288312
rect 0 287240 800 287360
rect 0 286152 800 286272
rect 0 285200 800 285320
rect 0 284112 800 284232
rect 0 283160 800 283280
rect 0 282072 800 282192
rect 0 281120 800 281240
rect 0 280032 800 280152
rect 0 279080 800 279200
rect 0 278128 800 278248
rect 0 277040 800 277160
rect 0 276088 800 276208
rect 0 275000 800 275120
rect 0 274048 800 274168
rect 0 272960 800 273080
rect 0 272008 800 272128
rect 0 270920 800 271040
rect 0 269968 800 270088
rect 0 268880 800 269000
rect 0 267928 800 268048
rect 0 266976 800 267096
rect 0 265888 800 266008
rect 0 264936 800 265056
rect 0 263848 800 263968
rect 0 262896 800 263016
rect 0 261808 800 261928
rect 0 260856 800 260976
rect 0 259768 800 259888
rect 0 258816 800 258936
rect 0 257728 800 257848
rect 0 256776 800 256896
rect 0 255824 800 255944
rect 0 254736 800 254856
rect 0 253784 800 253904
rect 0 252696 800 252816
rect 0 251744 800 251864
rect 0 250656 800 250776
rect 0 249704 800 249824
rect 0 248616 800 248736
rect 0 247664 800 247784
rect 0 246712 800 246832
rect 0 245624 800 245744
rect 0 244672 800 244792
rect 0 243584 800 243704
rect 0 242632 800 242752
rect 0 241544 800 241664
rect 0 240592 800 240712
rect 0 239504 800 239624
rect 0 238552 800 238672
rect 0 237464 800 237584
rect 0 236512 800 236632
rect 0 235560 800 235680
rect 0 234472 800 234592
rect 0 233520 800 233640
rect 0 232432 800 232552
rect 0 231480 800 231600
rect 0 230392 800 230512
rect 0 229440 800 229560
rect 0 228352 800 228472
rect 0 227400 800 227520
rect 0 226312 800 226432
rect 0 225360 800 225480
rect 0 224408 800 224528
rect 0 223320 800 223440
rect 0 222368 800 222488
rect 0 221280 800 221400
rect 0 220328 800 220448
rect 0 219240 800 219360
rect 0 218288 800 218408
rect 0 217200 800 217320
rect 0 216248 800 216368
rect 0 215160 800 215280
rect 0 214208 800 214328
rect 0 213256 800 213376
rect 0 212168 800 212288
rect 0 211216 800 211336
rect 0 210128 800 210248
rect 0 209176 800 209296
rect 0 208088 800 208208
rect 0 207136 800 207256
rect 0 206048 800 206168
rect 0 205096 800 205216
rect 0 204008 800 204128
rect 0 203056 800 203176
rect 0 202104 800 202224
rect 0 201016 800 201136
rect 0 200064 800 200184
rect 0 198976 800 199096
rect 0 198024 800 198144
rect 0 196936 800 197056
rect 0 195984 800 196104
rect 0 194896 800 195016
rect 0 193944 800 194064
rect 0 192992 800 193112
rect 0 191904 800 192024
rect 0 190952 800 191072
rect 0 189864 800 189984
rect 0 188912 800 189032
rect 0 187824 800 187944
rect 0 186872 800 186992
rect 0 185784 800 185904
rect 0 184832 800 184952
rect 0 183744 800 183864
rect 0 182792 800 182912
rect 0 181840 800 181960
rect 0 180752 800 180872
rect 0 179800 800 179920
rect 0 178712 800 178832
rect 0 177760 800 177880
rect 0 176672 800 176792
rect 0 175720 800 175840
rect 0 174632 800 174752
rect 0 173680 800 173800
rect 0 172592 800 172712
rect 0 171640 800 171760
rect 0 170688 800 170808
rect 0 169600 800 169720
rect 0 168648 800 168768
rect 0 167560 800 167680
rect 0 166608 800 166728
rect 0 165520 800 165640
rect 0 164568 800 164688
rect 0 163480 800 163600
rect 0 162528 800 162648
rect 0 161440 800 161560
rect 0 160488 800 160608
rect 0 159536 800 159656
rect 0 158448 800 158568
rect 0 157496 800 157616
rect 0 156408 800 156528
rect 0 155456 800 155576
rect 0 154368 800 154488
rect 0 153416 800 153536
rect 0 152328 800 152448
rect 0 151376 800 151496
rect 0 150424 800 150544
rect 0 149336 800 149456
rect 0 148384 800 148504
rect 0 147296 800 147416
rect 0 146344 800 146464
rect 0 145256 800 145376
rect 0 144304 800 144424
rect 0 143216 800 143336
rect 0 142264 800 142384
rect 0 141176 800 141296
rect 0 140224 800 140344
rect 0 139272 800 139392
rect 0 138184 800 138304
rect 0 137232 800 137352
rect 0 136144 800 136264
rect 0 135192 800 135312
rect 0 134104 800 134224
rect 0 133152 800 133272
rect 0 132064 800 132184
rect 0 131112 800 131232
rect 0 130024 800 130144
rect 0 129072 800 129192
rect 0 128120 800 128240
rect 0 127032 800 127152
rect 0 126080 800 126200
rect 0 124992 800 125112
rect 0 124040 800 124160
rect 0 122952 800 123072
rect 0 122000 800 122120
rect 0 120912 800 121032
rect 0 119960 800 120080
rect 0 118872 800 118992
rect 0 117920 800 118040
rect 0 116968 800 117088
rect 0 115880 800 116000
rect 0 114928 800 115048
rect 0 113840 800 113960
rect 0 112888 800 113008
rect 0 111800 800 111920
rect 0 110848 800 110968
rect 0 109760 800 109880
rect 0 108808 800 108928
rect 0 107720 800 107840
rect 0 106768 800 106888
rect 0 105816 800 105936
rect 0 104728 800 104848
rect 0 103776 800 103896
rect 0 102688 800 102808
rect 0 101736 800 101856
rect 0 100648 800 100768
rect 0 99696 800 99816
rect 0 98608 800 98728
rect 0 97656 800 97776
rect 0 96704 800 96824
rect 0 95616 800 95736
rect 0 94664 800 94784
rect 0 93576 800 93696
rect 0 92624 800 92744
rect 0 91536 800 91656
rect 0 90584 800 90704
rect 0 89496 800 89616
rect 0 88544 800 88664
rect 0 87456 800 87576
rect 0 86504 800 86624
rect 0 85552 800 85672
rect 0 84464 800 84584
rect 0 83512 800 83632
rect 0 82424 800 82544
rect 0 81472 800 81592
rect 0 80384 800 80504
rect 0 79432 800 79552
rect 0 78344 800 78464
rect 0 77392 800 77512
rect 0 76304 800 76424
rect 0 75352 800 75472
rect 0 74400 800 74520
rect 0 73312 800 73432
rect 0 72360 800 72480
rect 0 71272 800 71392
rect 0 70320 800 70440
rect 0 69232 800 69352
rect 0 68280 800 68400
rect 0 67192 800 67312
rect 0 66240 800 66360
rect 0 65152 800 65272
rect 0 64200 800 64320
rect 0 63248 800 63368
rect 0 62160 800 62280
rect 0 61208 800 61328
rect 0 60120 800 60240
rect 0 59168 800 59288
rect 0 58080 800 58200
rect 0 57128 800 57248
rect 0 56040 800 56160
rect 0 55088 800 55208
rect 0 54000 800 54120
rect 0 53048 800 53168
rect 0 52096 800 52216
rect 0 51008 800 51128
rect 0 50056 800 50176
rect 0 48968 800 49088
rect 0 48016 800 48136
rect 0 46928 800 47048
rect 0 45976 800 46096
rect 0 44888 800 45008
rect 0 43936 800 44056
rect 0 42984 800 43104
rect 0 41896 800 42016
rect 0 40944 800 41064
rect 0 39856 800 39976
rect 0 38904 800 39024
rect 0 37816 800 37936
rect 0 36864 800 36984
rect 0 35776 800 35896
rect 0 34824 800 34944
rect 0 33736 800 33856
rect 0 32784 800 32904
rect 0 31832 800 31952
rect 0 30744 800 30864
rect 0 29792 800 29912
rect 0 28704 800 28824
rect 0 27752 800 27872
rect 0 26664 800 26784
rect 0 25712 800 25832
rect 0 24624 800 24744
rect 0 23672 800 23792
rect 0 22584 800 22704
rect 0 21632 800 21752
rect 0 20680 800 20800
rect 0 19592 800 19712
rect 0 18640 800 18760
rect 0 17552 800 17672
rect 0 16600 800 16720
rect 0 15512 800 15632
rect 0 14560 800 14680
rect 0 13472 800 13592
rect 0 12520 800 12640
rect 0 11432 800 11552
rect 0 10480 800 10600
rect 0 9528 800 9648
rect 0 8440 800 8560
rect 0 7488 800 7608
rect 0 6400 800 6520
rect 0 5448 800 5568
rect 0 4360 800 4480
rect 0 3408 800 3528
rect 0 2320 800 2440
rect 0 1368 800 1488
rect 0 416 800 536
<< obsm3 >>
rect 880 299264 296368 299437
rect 800 298592 296368 299264
rect 880 298312 296368 298592
rect 800 297504 296368 298312
rect 880 297224 296368 297504
rect 800 296552 296368 297224
rect 880 296272 296368 296552
rect 800 295464 296368 296272
rect 880 295184 296368 295464
rect 800 294512 296368 295184
rect 880 294232 296368 294512
rect 800 293424 296368 294232
rect 880 293144 296368 293424
rect 800 292472 296368 293144
rect 880 292192 296368 292472
rect 800 291384 296368 292192
rect 880 291104 296368 291384
rect 800 290432 296368 291104
rect 880 290152 296368 290432
rect 800 289480 296368 290152
rect 880 289200 296368 289480
rect 800 288392 296368 289200
rect 880 288112 296368 288392
rect 800 287440 296368 288112
rect 880 287160 296368 287440
rect 800 286352 296368 287160
rect 880 286072 296368 286352
rect 800 285400 296368 286072
rect 880 285120 296368 285400
rect 800 284312 296368 285120
rect 880 284032 296368 284312
rect 800 283360 296368 284032
rect 880 283080 296368 283360
rect 800 282272 296368 283080
rect 880 281992 296368 282272
rect 800 281320 296368 281992
rect 880 281040 296368 281320
rect 800 280232 296368 281040
rect 880 279952 296368 280232
rect 800 279280 296368 279952
rect 880 279000 296368 279280
rect 800 278328 296368 279000
rect 880 278048 296368 278328
rect 800 277240 296368 278048
rect 880 276960 296368 277240
rect 800 276288 296368 276960
rect 880 276008 296368 276288
rect 800 275200 296368 276008
rect 880 274920 296368 275200
rect 800 274248 296368 274920
rect 880 273968 296368 274248
rect 800 273160 296368 273968
rect 880 272880 296368 273160
rect 800 272208 296368 272880
rect 880 271928 296368 272208
rect 800 271120 296368 271928
rect 880 270840 296368 271120
rect 800 270168 296368 270840
rect 880 269888 296368 270168
rect 800 269080 296368 269888
rect 880 268800 296368 269080
rect 800 268128 296368 268800
rect 880 267848 296368 268128
rect 800 267176 296368 267848
rect 880 266896 296368 267176
rect 800 266088 296368 266896
rect 880 265808 296368 266088
rect 800 265136 296368 265808
rect 880 264856 296368 265136
rect 800 264048 296368 264856
rect 880 263768 296368 264048
rect 800 263096 296368 263768
rect 880 262816 296368 263096
rect 800 262008 296368 262816
rect 880 261728 296368 262008
rect 800 261056 296368 261728
rect 880 260776 296368 261056
rect 800 259968 296368 260776
rect 880 259688 296368 259968
rect 800 259016 296368 259688
rect 880 258736 296368 259016
rect 800 257928 296368 258736
rect 880 257648 296368 257928
rect 800 256976 296368 257648
rect 880 256696 296368 256976
rect 800 256024 296368 256696
rect 880 255744 296368 256024
rect 800 254936 296368 255744
rect 880 254656 296368 254936
rect 800 253984 296368 254656
rect 880 253704 296368 253984
rect 800 252896 296368 253704
rect 880 252616 296368 252896
rect 800 251944 296368 252616
rect 880 251664 296368 251944
rect 800 250856 296368 251664
rect 880 250576 296368 250856
rect 800 249904 296368 250576
rect 880 249624 296368 249904
rect 800 248816 296368 249624
rect 880 248536 296368 248816
rect 800 247864 296368 248536
rect 880 247584 296368 247864
rect 800 246912 296368 247584
rect 880 246632 296368 246912
rect 800 245824 296368 246632
rect 880 245544 296368 245824
rect 800 244872 296368 245544
rect 880 244592 296368 244872
rect 800 243784 296368 244592
rect 880 243504 296368 243784
rect 800 242832 296368 243504
rect 880 242552 296368 242832
rect 800 241744 296368 242552
rect 880 241464 296368 241744
rect 800 240792 296368 241464
rect 880 240512 296368 240792
rect 800 239704 296368 240512
rect 880 239424 296368 239704
rect 800 238752 296368 239424
rect 880 238472 296368 238752
rect 800 237664 296368 238472
rect 880 237384 296368 237664
rect 800 236712 296368 237384
rect 880 236432 296368 236712
rect 800 235760 296368 236432
rect 880 235480 296368 235760
rect 800 234672 296368 235480
rect 880 234392 296368 234672
rect 800 233720 296368 234392
rect 880 233440 296368 233720
rect 800 232632 296368 233440
rect 880 232352 296368 232632
rect 800 231680 296368 232352
rect 880 231400 296368 231680
rect 800 230592 296368 231400
rect 880 230312 296368 230592
rect 800 229640 296368 230312
rect 880 229360 296368 229640
rect 800 228552 296368 229360
rect 880 228272 296368 228552
rect 800 227600 296368 228272
rect 880 227320 296368 227600
rect 800 226512 296368 227320
rect 880 226232 296368 226512
rect 800 225560 296368 226232
rect 880 225280 296368 225560
rect 800 224608 296368 225280
rect 880 224328 296368 224608
rect 800 223520 296368 224328
rect 880 223240 296368 223520
rect 800 222568 296368 223240
rect 880 222288 296368 222568
rect 800 221480 296368 222288
rect 880 221200 296368 221480
rect 800 220528 296368 221200
rect 880 220248 296368 220528
rect 800 219440 296368 220248
rect 880 219160 296368 219440
rect 800 218488 296368 219160
rect 880 218208 296368 218488
rect 800 217400 296368 218208
rect 880 217120 296368 217400
rect 800 216448 296368 217120
rect 880 216168 296368 216448
rect 800 215360 296368 216168
rect 880 215080 296368 215360
rect 800 214408 296368 215080
rect 880 214128 296368 214408
rect 800 213456 296368 214128
rect 880 213176 296368 213456
rect 800 212368 296368 213176
rect 880 212088 296368 212368
rect 800 211416 296368 212088
rect 880 211136 296368 211416
rect 800 210328 296368 211136
rect 880 210048 296368 210328
rect 800 209376 296368 210048
rect 880 209096 296368 209376
rect 800 208288 296368 209096
rect 880 208008 296368 208288
rect 800 207336 296368 208008
rect 880 207056 296368 207336
rect 800 206248 296368 207056
rect 880 205968 296368 206248
rect 800 205296 296368 205968
rect 880 205016 296368 205296
rect 800 204208 296368 205016
rect 880 203928 296368 204208
rect 800 203256 296368 203928
rect 880 202976 296368 203256
rect 800 202304 296368 202976
rect 880 202024 296368 202304
rect 800 201216 296368 202024
rect 880 200936 296368 201216
rect 800 200264 296368 200936
rect 880 199984 296368 200264
rect 800 199176 296368 199984
rect 880 198896 296368 199176
rect 800 198224 296368 198896
rect 880 197944 296368 198224
rect 800 197136 296368 197944
rect 880 196856 296368 197136
rect 800 196184 296368 196856
rect 880 195904 296368 196184
rect 800 195096 296368 195904
rect 880 194816 296368 195096
rect 800 194144 296368 194816
rect 880 193864 296368 194144
rect 800 193192 296368 193864
rect 880 192912 296368 193192
rect 800 192104 296368 192912
rect 880 191824 296368 192104
rect 800 191152 296368 191824
rect 880 190872 296368 191152
rect 800 190064 296368 190872
rect 880 189784 296368 190064
rect 800 189112 296368 189784
rect 880 188832 296368 189112
rect 800 188024 296368 188832
rect 880 187744 296368 188024
rect 800 187072 296368 187744
rect 880 186792 296368 187072
rect 800 185984 296368 186792
rect 880 185704 296368 185984
rect 800 185032 296368 185704
rect 880 184752 296368 185032
rect 800 183944 296368 184752
rect 880 183664 296368 183944
rect 800 182992 296368 183664
rect 880 182712 296368 182992
rect 800 182040 296368 182712
rect 880 181760 296368 182040
rect 800 180952 296368 181760
rect 880 180672 296368 180952
rect 800 180000 296368 180672
rect 880 179720 296368 180000
rect 800 178912 296368 179720
rect 880 178632 296368 178912
rect 800 177960 296368 178632
rect 880 177680 296368 177960
rect 800 176872 296368 177680
rect 880 176592 296368 176872
rect 800 175920 296368 176592
rect 880 175640 296368 175920
rect 800 174832 296368 175640
rect 880 174552 296368 174832
rect 800 173880 296368 174552
rect 880 173600 296368 173880
rect 800 172792 296368 173600
rect 880 172512 296368 172792
rect 800 171840 296368 172512
rect 880 171560 296368 171840
rect 800 170888 296368 171560
rect 880 170608 296368 170888
rect 800 169800 296368 170608
rect 880 169520 296368 169800
rect 800 168848 296368 169520
rect 880 168568 296368 168848
rect 800 167760 296368 168568
rect 880 167480 296368 167760
rect 800 166808 296368 167480
rect 880 166528 296368 166808
rect 800 165720 296368 166528
rect 880 165440 296368 165720
rect 800 164768 296368 165440
rect 880 164488 296368 164768
rect 800 163680 296368 164488
rect 880 163400 296368 163680
rect 800 162728 296368 163400
rect 880 162448 296368 162728
rect 800 161640 296368 162448
rect 880 161360 296368 161640
rect 800 160688 296368 161360
rect 880 160408 296368 160688
rect 800 159736 296368 160408
rect 880 159456 296368 159736
rect 800 158648 296368 159456
rect 880 158368 296368 158648
rect 800 157696 296368 158368
rect 880 157416 296368 157696
rect 800 156608 296368 157416
rect 880 156328 296368 156608
rect 800 155656 296368 156328
rect 880 155376 296368 155656
rect 800 154568 296368 155376
rect 880 154288 296368 154568
rect 800 153616 296368 154288
rect 880 153336 296368 153616
rect 800 152528 296368 153336
rect 880 152248 296368 152528
rect 800 151576 296368 152248
rect 880 151296 296368 151576
rect 800 150624 296368 151296
rect 880 150344 296368 150624
rect 800 149536 296368 150344
rect 880 149256 296368 149536
rect 800 148584 296368 149256
rect 880 148304 296368 148584
rect 800 147496 296368 148304
rect 880 147216 296368 147496
rect 800 146544 296368 147216
rect 880 146264 296368 146544
rect 800 145456 296368 146264
rect 880 145176 296368 145456
rect 800 144504 296368 145176
rect 880 144224 296368 144504
rect 800 143416 296368 144224
rect 880 143136 296368 143416
rect 800 142464 296368 143136
rect 880 142184 296368 142464
rect 800 141376 296368 142184
rect 880 141096 296368 141376
rect 800 140424 296368 141096
rect 880 140144 296368 140424
rect 800 139472 296368 140144
rect 880 139192 296368 139472
rect 800 138384 296368 139192
rect 880 138104 296368 138384
rect 800 137432 296368 138104
rect 880 137152 296368 137432
rect 800 136344 296368 137152
rect 880 136064 296368 136344
rect 800 135392 296368 136064
rect 880 135112 296368 135392
rect 800 134304 296368 135112
rect 880 134024 296368 134304
rect 800 133352 296368 134024
rect 880 133072 296368 133352
rect 800 132264 296368 133072
rect 880 131984 296368 132264
rect 800 131312 296368 131984
rect 880 131032 296368 131312
rect 800 130224 296368 131032
rect 880 129944 296368 130224
rect 800 129272 296368 129944
rect 880 128992 296368 129272
rect 800 128320 296368 128992
rect 880 128040 296368 128320
rect 800 127232 296368 128040
rect 880 126952 296368 127232
rect 800 126280 296368 126952
rect 880 126000 296368 126280
rect 800 125192 296368 126000
rect 880 124912 296368 125192
rect 800 124240 296368 124912
rect 880 123960 296368 124240
rect 800 123152 296368 123960
rect 880 122872 296368 123152
rect 800 122200 296368 122872
rect 880 121920 296368 122200
rect 800 121112 296368 121920
rect 880 120832 296368 121112
rect 800 120160 296368 120832
rect 880 119880 296368 120160
rect 800 119072 296368 119880
rect 880 118792 296368 119072
rect 800 118120 296368 118792
rect 880 117840 296368 118120
rect 800 117168 296368 117840
rect 880 116888 296368 117168
rect 800 116080 296368 116888
rect 880 115800 296368 116080
rect 800 115128 296368 115800
rect 880 114848 296368 115128
rect 800 114040 296368 114848
rect 880 113760 296368 114040
rect 800 113088 296368 113760
rect 880 112808 296368 113088
rect 800 112000 296368 112808
rect 880 111720 296368 112000
rect 800 111048 296368 111720
rect 880 110768 296368 111048
rect 800 109960 296368 110768
rect 880 109680 296368 109960
rect 800 109008 296368 109680
rect 880 108728 296368 109008
rect 800 107920 296368 108728
rect 880 107640 296368 107920
rect 800 106968 296368 107640
rect 880 106688 296368 106968
rect 800 106016 296368 106688
rect 880 105736 296368 106016
rect 800 104928 296368 105736
rect 880 104648 296368 104928
rect 800 103976 296368 104648
rect 880 103696 296368 103976
rect 800 102888 296368 103696
rect 880 102608 296368 102888
rect 800 101936 296368 102608
rect 880 101656 296368 101936
rect 800 100848 296368 101656
rect 880 100568 296368 100848
rect 800 99896 296368 100568
rect 880 99616 296368 99896
rect 800 98808 296368 99616
rect 880 98528 296368 98808
rect 800 97856 296368 98528
rect 880 97576 296368 97856
rect 800 96904 296368 97576
rect 880 96624 296368 96904
rect 800 95816 296368 96624
rect 880 95536 296368 95816
rect 800 94864 296368 95536
rect 880 94584 296368 94864
rect 800 93776 296368 94584
rect 880 93496 296368 93776
rect 800 92824 296368 93496
rect 880 92544 296368 92824
rect 800 91736 296368 92544
rect 880 91456 296368 91736
rect 800 90784 296368 91456
rect 880 90504 296368 90784
rect 800 89696 296368 90504
rect 880 89416 296368 89696
rect 800 88744 296368 89416
rect 880 88464 296368 88744
rect 800 87656 296368 88464
rect 880 87376 296368 87656
rect 800 86704 296368 87376
rect 880 86424 296368 86704
rect 800 85752 296368 86424
rect 880 85472 296368 85752
rect 800 84664 296368 85472
rect 880 84384 296368 84664
rect 800 83712 296368 84384
rect 880 83432 296368 83712
rect 800 82624 296368 83432
rect 880 82344 296368 82624
rect 800 81672 296368 82344
rect 880 81392 296368 81672
rect 800 80584 296368 81392
rect 880 80304 296368 80584
rect 800 79632 296368 80304
rect 880 79352 296368 79632
rect 800 78544 296368 79352
rect 880 78264 296368 78544
rect 800 77592 296368 78264
rect 880 77312 296368 77592
rect 800 76504 296368 77312
rect 880 76224 296368 76504
rect 800 75552 296368 76224
rect 880 75272 296368 75552
rect 800 74600 296368 75272
rect 880 74320 296368 74600
rect 800 73512 296368 74320
rect 880 73232 296368 73512
rect 800 72560 296368 73232
rect 880 72280 296368 72560
rect 800 71472 296368 72280
rect 880 71192 296368 71472
rect 800 70520 296368 71192
rect 880 70240 296368 70520
rect 800 69432 296368 70240
rect 880 69152 296368 69432
rect 800 68480 296368 69152
rect 880 68200 296368 68480
rect 800 67392 296368 68200
rect 880 67112 296368 67392
rect 800 66440 296368 67112
rect 880 66160 296368 66440
rect 800 65352 296368 66160
rect 880 65072 296368 65352
rect 800 64400 296368 65072
rect 880 64120 296368 64400
rect 800 63448 296368 64120
rect 880 63168 296368 63448
rect 800 62360 296368 63168
rect 880 62080 296368 62360
rect 800 61408 296368 62080
rect 880 61128 296368 61408
rect 800 60320 296368 61128
rect 880 60040 296368 60320
rect 800 59368 296368 60040
rect 880 59088 296368 59368
rect 800 58280 296368 59088
rect 880 58000 296368 58280
rect 800 57328 296368 58000
rect 880 57048 296368 57328
rect 800 56240 296368 57048
rect 880 55960 296368 56240
rect 800 55288 296368 55960
rect 880 55008 296368 55288
rect 800 54200 296368 55008
rect 880 53920 296368 54200
rect 800 53248 296368 53920
rect 880 52968 296368 53248
rect 800 52296 296368 52968
rect 880 52016 296368 52296
rect 800 51208 296368 52016
rect 880 50928 296368 51208
rect 800 50256 296368 50928
rect 880 49976 296368 50256
rect 800 49168 296368 49976
rect 880 48888 296368 49168
rect 800 48216 296368 48888
rect 880 47936 296368 48216
rect 800 47128 296368 47936
rect 880 46848 296368 47128
rect 800 46176 296368 46848
rect 880 45896 296368 46176
rect 800 45088 296368 45896
rect 880 44808 296368 45088
rect 800 44136 296368 44808
rect 880 43856 296368 44136
rect 800 43184 296368 43856
rect 880 42904 296368 43184
rect 800 42096 296368 42904
rect 880 41816 296368 42096
rect 800 41144 296368 41816
rect 880 40864 296368 41144
rect 800 40056 296368 40864
rect 880 39776 296368 40056
rect 800 39104 296368 39776
rect 880 38824 296368 39104
rect 800 38016 296368 38824
rect 880 37736 296368 38016
rect 800 37064 296368 37736
rect 880 36784 296368 37064
rect 800 35976 296368 36784
rect 880 35696 296368 35976
rect 800 35024 296368 35696
rect 880 34744 296368 35024
rect 800 33936 296368 34744
rect 880 33656 296368 33936
rect 800 32984 296368 33656
rect 880 32704 296368 32984
rect 800 32032 296368 32704
rect 880 31752 296368 32032
rect 800 30944 296368 31752
rect 880 30664 296368 30944
rect 800 29992 296368 30664
rect 880 29712 296368 29992
rect 800 28904 296368 29712
rect 880 28624 296368 28904
rect 800 27952 296368 28624
rect 880 27672 296368 27952
rect 800 26864 296368 27672
rect 880 26584 296368 26864
rect 800 25912 296368 26584
rect 880 25632 296368 25912
rect 800 24824 296368 25632
rect 880 24544 296368 24824
rect 800 23872 296368 24544
rect 880 23592 296368 23872
rect 800 22784 296368 23592
rect 880 22504 296368 22784
rect 800 21832 296368 22504
rect 880 21552 296368 21832
rect 800 20880 296368 21552
rect 880 20600 296368 20880
rect 800 19792 296368 20600
rect 880 19512 296368 19792
rect 800 18840 296368 19512
rect 880 18560 296368 18840
rect 800 17752 296368 18560
rect 880 17472 296368 17752
rect 800 16800 296368 17472
rect 880 16520 296368 16800
rect 800 15712 296368 16520
rect 880 15432 296368 15712
rect 800 14760 296368 15432
rect 880 14480 296368 14760
rect 800 13672 296368 14480
rect 880 13392 296368 13672
rect 800 12720 296368 13392
rect 880 12440 296368 12720
rect 800 11632 296368 12440
rect 880 11352 296368 11632
rect 800 10680 296368 11352
rect 880 10400 296368 10680
rect 800 9728 296368 10400
rect 880 9448 296368 9728
rect 800 8640 296368 9448
rect 880 8360 296368 8640
rect 800 7688 296368 8360
rect 880 7408 296368 7688
rect 800 6600 296368 7408
rect 880 6320 296368 6600
rect 800 5648 296368 6320
rect 880 5368 296368 5648
rect 800 4560 296368 5368
rect 880 4280 296368 4560
rect 800 3608 296368 4280
rect 880 3328 296368 3608
rect 800 2520 296368 3328
rect 880 2240 296368 2520
rect 800 1568 296368 2240
rect 880 1288 296368 1568
rect 800 616 296368 1288
rect 880 443 296368 616
<< metal4 >>
rect 4208 2128 4528 297616
rect 19568 2128 19888 297616
rect 34928 2128 35248 297616
rect 50288 2128 50608 297616
rect 65648 2128 65968 297616
rect 81008 2128 81328 297616
rect 96368 2128 96688 297616
rect 111728 2128 112048 297616
rect 127088 2128 127408 297616
rect 142448 2128 142768 297616
rect 157808 2128 158128 297616
rect 173168 2128 173488 297616
rect 188528 2128 188848 297616
rect 203888 2128 204208 297616
rect 219248 2128 219568 297616
rect 234608 2128 234928 297616
rect 249968 2128 250288 297616
rect 265328 2128 265648 297616
rect 280688 2128 281008 297616
rect 296048 2128 296368 297616
<< obsm4 >>
rect 979 2619 4128 296853
rect 4608 2619 19488 296853
rect 19968 2619 34848 296853
rect 35328 2619 50208 296853
rect 50688 2619 65568 296853
rect 66048 2619 80928 296853
rect 81408 2619 96288 296853
rect 96768 2619 111648 296853
rect 112128 2619 127008 296853
rect 127488 2619 142368 296853
rect 142848 2619 157728 296853
rect 158208 2619 173088 296853
rect 173568 2619 178053 296853
<< labels >>
rlabel metal3 s 0 134104 800 134224 6 bb_addr0[0]
port 1 nsew signal output
rlabel metal3 s 0 188912 800 189032 6 bb_addr0[10]
port 2 nsew signal output
rlabel metal3 s 0 193944 800 194064 6 bb_addr0[11]
port 3 nsew signal output
rlabel metal3 s 0 198976 800 199096 6 bb_addr0[12]
port 4 nsew signal output
rlabel metal3 s 0 204008 800 204128 6 bb_addr0[13]
port 5 nsew signal output
rlabel metal3 s 0 209176 800 209296 6 bb_addr0[14]
port 6 nsew signal output
rlabel metal3 s 0 214208 800 214328 6 bb_addr0[15]
port 7 nsew signal output
rlabel metal3 s 0 219240 800 219360 6 bb_addr0[16]
port 8 nsew signal output
rlabel metal3 s 0 224408 800 224528 6 bb_addr0[17]
port 9 nsew signal output
rlabel metal3 s 0 229440 800 229560 6 bb_addr0[18]
port 10 nsew signal output
rlabel metal3 s 0 234472 800 234592 6 bb_addr0[19]
port 11 nsew signal output
rlabel metal3 s 0 140224 800 140344 6 bb_addr0[1]
port 12 nsew signal output
rlabel metal3 s 0 239504 800 239624 6 bb_addr0[20]
port 13 nsew signal output
rlabel metal3 s 0 244672 800 244792 6 bb_addr0[21]
port 14 nsew signal output
rlabel metal3 s 0 249704 800 249824 6 bb_addr0[22]
port 15 nsew signal output
rlabel metal3 s 0 254736 800 254856 6 bb_addr0[23]
port 16 nsew signal output
rlabel metal3 s 0 259768 800 259888 6 bb_addr0[24]
port 17 nsew signal output
rlabel metal3 s 0 264936 800 265056 6 bb_addr0[25]
port 18 nsew signal output
rlabel metal3 s 0 269968 800 270088 6 bb_addr0[26]
port 19 nsew signal output
rlabel metal3 s 0 275000 800 275120 6 bb_addr0[27]
port 20 nsew signal output
rlabel metal3 s 0 280032 800 280152 6 bb_addr0[28]
port 21 nsew signal output
rlabel metal3 s 0 285200 800 285320 6 bb_addr0[29]
port 22 nsew signal output
rlabel metal3 s 0 146344 800 146464 6 bb_addr0[2]
port 23 nsew signal output
rlabel metal3 s 0 290232 800 290352 6 bb_addr0[30]
port 24 nsew signal output
rlabel metal3 s 0 295264 800 295384 6 bb_addr0[31]
port 25 nsew signal output
rlabel metal3 s 0 152328 800 152448 6 bb_addr0[3]
port 26 nsew signal output
rlabel metal3 s 0 158448 800 158568 6 bb_addr0[4]
port 27 nsew signal output
rlabel metal3 s 0 163480 800 163600 6 bb_addr0[5]
port 28 nsew signal output
rlabel metal3 s 0 168648 800 168768 6 bb_addr0[6]
port 29 nsew signal output
rlabel metal3 s 0 173680 800 173800 6 bb_addr0[7]
port 30 nsew signal output
rlabel metal3 s 0 178712 800 178832 6 bb_addr0[8]
port 31 nsew signal output
rlabel metal3 s 0 183744 800 183864 6 bb_addr0[9]
port 32 nsew signal output
rlabel metal3 s 0 135192 800 135312 6 bb_addr1[0]
port 33 nsew signal output
rlabel metal3 s 0 189864 800 189984 6 bb_addr1[10]
port 34 nsew signal output
rlabel metal3 s 0 194896 800 195016 6 bb_addr1[11]
port 35 nsew signal output
rlabel metal3 s 0 200064 800 200184 6 bb_addr1[12]
port 36 nsew signal output
rlabel metal3 s 0 205096 800 205216 6 bb_addr1[13]
port 37 nsew signal output
rlabel metal3 s 0 210128 800 210248 6 bb_addr1[14]
port 38 nsew signal output
rlabel metal3 s 0 215160 800 215280 6 bb_addr1[15]
port 39 nsew signal output
rlabel metal3 s 0 220328 800 220448 6 bb_addr1[16]
port 40 nsew signal output
rlabel metal3 s 0 225360 800 225480 6 bb_addr1[17]
port 41 nsew signal output
rlabel metal3 s 0 230392 800 230512 6 bb_addr1[18]
port 42 nsew signal output
rlabel metal3 s 0 235560 800 235680 6 bb_addr1[19]
port 43 nsew signal output
rlabel metal3 s 0 141176 800 141296 6 bb_addr1[1]
port 44 nsew signal output
rlabel metal3 s 0 240592 800 240712 6 bb_addr1[20]
port 45 nsew signal output
rlabel metal3 s 0 245624 800 245744 6 bb_addr1[21]
port 46 nsew signal output
rlabel metal3 s 0 250656 800 250776 6 bb_addr1[22]
port 47 nsew signal output
rlabel metal3 s 0 255824 800 255944 6 bb_addr1[23]
port 48 nsew signal output
rlabel metal3 s 0 260856 800 260976 6 bb_addr1[24]
port 49 nsew signal output
rlabel metal3 s 0 265888 800 266008 6 bb_addr1[25]
port 50 nsew signal output
rlabel metal3 s 0 270920 800 271040 6 bb_addr1[26]
port 51 nsew signal output
rlabel metal3 s 0 276088 800 276208 6 bb_addr1[27]
port 52 nsew signal output
rlabel metal3 s 0 281120 800 281240 6 bb_addr1[28]
port 53 nsew signal output
rlabel metal3 s 0 286152 800 286272 6 bb_addr1[29]
port 54 nsew signal output
rlabel metal3 s 0 147296 800 147416 6 bb_addr1[2]
port 55 nsew signal output
rlabel metal3 s 0 291184 800 291304 6 bb_addr1[30]
port 56 nsew signal output
rlabel metal3 s 0 296352 800 296472 6 bb_addr1[31]
port 57 nsew signal output
rlabel metal3 s 0 153416 800 153536 6 bb_addr1[3]
port 58 nsew signal output
rlabel metal3 s 0 159536 800 159656 6 bb_addr1[4]
port 59 nsew signal output
rlabel metal3 s 0 164568 800 164688 6 bb_addr1[5]
port 60 nsew signal output
rlabel metal3 s 0 169600 800 169720 6 bb_addr1[6]
port 61 nsew signal output
rlabel metal3 s 0 174632 800 174752 6 bb_addr1[7]
port 62 nsew signal output
rlabel metal3 s 0 179800 800 179920 6 bb_addr1[8]
port 63 nsew signal output
rlabel metal3 s 0 184832 800 184952 6 bb_addr1[9]
port 64 nsew signal output
rlabel metal3 s 0 131112 800 131232 6 bb_csb0
port 65 nsew signal output
rlabel metal3 s 0 132064 800 132184 6 bb_csb1
port 66 nsew signal output
rlabel metal3 s 0 136144 800 136264 6 bb_din0[0]
port 67 nsew signal output
rlabel metal3 s 0 190952 800 191072 6 bb_din0[10]
port 68 nsew signal output
rlabel metal3 s 0 195984 800 196104 6 bb_din0[11]
port 69 nsew signal output
rlabel metal3 s 0 201016 800 201136 6 bb_din0[12]
port 70 nsew signal output
rlabel metal3 s 0 206048 800 206168 6 bb_din0[13]
port 71 nsew signal output
rlabel metal3 s 0 211216 800 211336 6 bb_din0[14]
port 72 nsew signal output
rlabel metal3 s 0 216248 800 216368 6 bb_din0[15]
port 73 nsew signal output
rlabel metal3 s 0 221280 800 221400 6 bb_din0[16]
port 74 nsew signal output
rlabel metal3 s 0 226312 800 226432 6 bb_din0[17]
port 75 nsew signal output
rlabel metal3 s 0 231480 800 231600 6 bb_din0[18]
port 76 nsew signal output
rlabel metal3 s 0 236512 800 236632 6 bb_din0[19]
port 77 nsew signal output
rlabel metal3 s 0 142264 800 142384 6 bb_din0[1]
port 78 nsew signal output
rlabel metal3 s 0 241544 800 241664 6 bb_din0[20]
port 79 nsew signal output
rlabel metal3 s 0 246712 800 246832 6 bb_din0[21]
port 80 nsew signal output
rlabel metal3 s 0 251744 800 251864 6 bb_din0[22]
port 81 nsew signal output
rlabel metal3 s 0 256776 800 256896 6 bb_din0[23]
port 82 nsew signal output
rlabel metal3 s 0 261808 800 261928 6 bb_din0[24]
port 83 nsew signal output
rlabel metal3 s 0 266976 800 267096 6 bb_din0[25]
port 84 nsew signal output
rlabel metal3 s 0 272008 800 272128 6 bb_din0[26]
port 85 nsew signal output
rlabel metal3 s 0 277040 800 277160 6 bb_din0[27]
port 86 nsew signal output
rlabel metal3 s 0 282072 800 282192 6 bb_din0[28]
port 87 nsew signal output
rlabel metal3 s 0 287240 800 287360 6 bb_din0[29]
port 88 nsew signal output
rlabel metal3 s 0 148384 800 148504 6 bb_din0[2]
port 89 nsew signal output
rlabel metal3 s 0 292272 800 292392 6 bb_din0[30]
port 90 nsew signal output
rlabel metal3 s 0 297304 800 297424 6 bb_din0[31]
port 91 nsew signal output
rlabel metal3 s 0 154368 800 154488 6 bb_din0[3]
port 92 nsew signal output
rlabel metal3 s 0 160488 800 160608 6 bb_din0[4]
port 93 nsew signal output
rlabel metal3 s 0 165520 800 165640 6 bb_din0[5]
port 94 nsew signal output
rlabel metal3 s 0 170688 800 170808 6 bb_din0[6]
port 95 nsew signal output
rlabel metal3 s 0 175720 800 175840 6 bb_din0[7]
port 96 nsew signal output
rlabel metal3 s 0 180752 800 180872 6 bb_din0[8]
port 97 nsew signal output
rlabel metal3 s 0 185784 800 185904 6 bb_din0[9]
port 98 nsew signal output
rlabel metal3 s 0 137232 800 137352 6 bb_dout0[0]
port 99 nsew signal input
rlabel metal3 s 0 191904 800 192024 6 bb_dout0[10]
port 100 nsew signal input
rlabel metal3 s 0 196936 800 197056 6 bb_dout0[11]
port 101 nsew signal input
rlabel metal3 s 0 202104 800 202224 6 bb_dout0[12]
port 102 nsew signal input
rlabel metal3 s 0 207136 800 207256 6 bb_dout0[13]
port 103 nsew signal input
rlabel metal3 s 0 212168 800 212288 6 bb_dout0[14]
port 104 nsew signal input
rlabel metal3 s 0 217200 800 217320 6 bb_dout0[15]
port 105 nsew signal input
rlabel metal3 s 0 222368 800 222488 6 bb_dout0[16]
port 106 nsew signal input
rlabel metal3 s 0 227400 800 227520 6 bb_dout0[17]
port 107 nsew signal input
rlabel metal3 s 0 232432 800 232552 6 bb_dout0[18]
port 108 nsew signal input
rlabel metal3 s 0 237464 800 237584 6 bb_dout0[19]
port 109 nsew signal input
rlabel metal3 s 0 143216 800 143336 6 bb_dout0[1]
port 110 nsew signal input
rlabel metal3 s 0 242632 800 242752 6 bb_dout0[20]
port 111 nsew signal input
rlabel metal3 s 0 247664 800 247784 6 bb_dout0[21]
port 112 nsew signal input
rlabel metal3 s 0 252696 800 252816 6 bb_dout0[22]
port 113 nsew signal input
rlabel metal3 s 0 257728 800 257848 6 bb_dout0[23]
port 114 nsew signal input
rlabel metal3 s 0 262896 800 263016 6 bb_dout0[24]
port 115 nsew signal input
rlabel metal3 s 0 267928 800 268048 6 bb_dout0[25]
port 116 nsew signal input
rlabel metal3 s 0 272960 800 273080 6 bb_dout0[26]
port 117 nsew signal input
rlabel metal3 s 0 278128 800 278248 6 bb_dout0[27]
port 118 nsew signal input
rlabel metal3 s 0 283160 800 283280 6 bb_dout0[28]
port 119 nsew signal input
rlabel metal3 s 0 288192 800 288312 6 bb_dout0[29]
port 120 nsew signal input
rlabel metal3 s 0 149336 800 149456 6 bb_dout0[2]
port 121 nsew signal input
rlabel metal3 s 0 293224 800 293344 6 bb_dout0[30]
port 122 nsew signal input
rlabel metal3 s 0 298392 800 298512 6 bb_dout0[31]
port 123 nsew signal input
rlabel metal3 s 0 155456 800 155576 6 bb_dout0[3]
port 124 nsew signal input
rlabel metal3 s 0 161440 800 161560 6 bb_dout0[4]
port 125 nsew signal input
rlabel metal3 s 0 166608 800 166728 6 bb_dout0[5]
port 126 nsew signal input
rlabel metal3 s 0 171640 800 171760 6 bb_dout0[6]
port 127 nsew signal input
rlabel metal3 s 0 176672 800 176792 6 bb_dout0[7]
port 128 nsew signal input
rlabel metal3 s 0 181840 800 181960 6 bb_dout0[8]
port 129 nsew signal input
rlabel metal3 s 0 186872 800 186992 6 bb_dout0[9]
port 130 nsew signal input
rlabel metal3 s 0 138184 800 138304 6 bb_dout1[0]
port 131 nsew signal input
rlabel metal3 s 0 192992 800 193112 6 bb_dout1[10]
port 132 nsew signal input
rlabel metal3 s 0 198024 800 198144 6 bb_dout1[11]
port 133 nsew signal input
rlabel metal3 s 0 203056 800 203176 6 bb_dout1[12]
port 134 nsew signal input
rlabel metal3 s 0 208088 800 208208 6 bb_dout1[13]
port 135 nsew signal input
rlabel metal3 s 0 213256 800 213376 6 bb_dout1[14]
port 136 nsew signal input
rlabel metal3 s 0 218288 800 218408 6 bb_dout1[15]
port 137 nsew signal input
rlabel metal3 s 0 223320 800 223440 6 bb_dout1[16]
port 138 nsew signal input
rlabel metal3 s 0 228352 800 228472 6 bb_dout1[17]
port 139 nsew signal input
rlabel metal3 s 0 233520 800 233640 6 bb_dout1[18]
port 140 nsew signal input
rlabel metal3 s 0 238552 800 238672 6 bb_dout1[19]
port 141 nsew signal input
rlabel metal3 s 0 144304 800 144424 6 bb_dout1[1]
port 142 nsew signal input
rlabel metal3 s 0 243584 800 243704 6 bb_dout1[20]
port 143 nsew signal input
rlabel metal3 s 0 248616 800 248736 6 bb_dout1[21]
port 144 nsew signal input
rlabel metal3 s 0 253784 800 253904 6 bb_dout1[22]
port 145 nsew signal input
rlabel metal3 s 0 258816 800 258936 6 bb_dout1[23]
port 146 nsew signal input
rlabel metal3 s 0 263848 800 263968 6 bb_dout1[24]
port 147 nsew signal input
rlabel metal3 s 0 268880 800 269000 6 bb_dout1[25]
port 148 nsew signal input
rlabel metal3 s 0 274048 800 274168 6 bb_dout1[26]
port 149 nsew signal input
rlabel metal3 s 0 279080 800 279200 6 bb_dout1[27]
port 150 nsew signal input
rlabel metal3 s 0 284112 800 284232 6 bb_dout1[28]
port 151 nsew signal input
rlabel metal3 s 0 289280 800 289400 6 bb_dout1[29]
port 152 nsew signal input
rlabel metal3 s 0 150424 800 150544 6 bb_dout1[2]
port 153 nsew signal input
rlabel metal3 s 0 294312 800 294432 6 bb_dout1[30]
port 154 nsew signal input
rlabel metal3 s 0 299344 800 299464 6 bb_dout1[31]
port 155 nsew signal input
rlabel metal3 s 0 156408 800 156528 6 bb_dout1[3]
port 156 nsew signal input
rlabel metal3 s 0 162528 800 162648 6 bb_dout1[4]
port 157 nsew signal input
rlabel metal3 s 0 167560 800 167680 6 bb_dout1[5]
port 158 nsew signal input
rlabel metal3 s 0 172592 800 172712 6 bb_dout1[6]
port 159 nsew signal input
rlabel metal3 s 0 177760 800 177880 6 bb_dout1[7]
port 160 nsew signal input
rlabel metal3 s 0 182792 800 182912 6 bb_dout1[8]
port 161 nsew signal input
rlabel metal3 s 0 187824 800 187944 6 bb_dout1[9]
port 162 nsew signal input
rlabel metal3 s 0 133152 800 133272 6 bb_web0
port 163 nsew signal output
rlabel metal3 s 0 139272 800 139392 6 bb_wmask0[0]
port 164 nsew signal output
rlabel metal3 s 0 145256 800 145376 6 bb_wmask0[1]
port 165 nsew signal output
rlabel metal3 s 0 151376 800 151496 6 bb_wmask0[2]
port 166 nsew signal output
rlabel metal3 s 0 157496 800 157616 6 bb_wmask0[3]
port 167 nsew signal output
rlabel metal2 s 1950 0 2006 800 6 clk_g
port 168 nsew signal input
rlabel metal2 s 17866 0 17922 800 6 io_gecerli
port 169 nsew signal output
rlabel metal2 s 21914 0 21970 800 6 io_oeb[0]
port 170 nsew signal output
rlabel metal2 s 101954 0 102010 800 6 io_oeb[10]
port 171 nsew signal output
rlabel metal2 s 109866 0 109922 800 6 io_oeb[11]
port 172 nsew signal output
rlabel metal2 s 117870 0 117926 800 6 io_oeb[12]
port 173 nsew signal output
rlabel metal2 s 125874 0 125930 800 6 io_oeb[13]
port 174 nsew signal output
rlabel metal2 s 133878 0 133934 800 6 io_oeb[14]
port 175 nsew signal output
rlabel metal2 s 141882 0 141938 800 6 io_oeb[15]
port 176 nsew signal output
rlabel metal2 s 149886 0 149942 800 6 io_oeb[16]
port 177 nsew signal output
rlabel metal2 s 157890 0 157946 800 6 io_oeb[17]
port 178 nsew signal output
rlabel metal2 s 165894 0 165950 800 6 io_oeb[18]
port 179 nsew signal output
rlabel metal2 s 173898 0 173954 800 6 io_oeb[19]
port 180 nsew signal output
rlabel metal2 s 29918 0 29974 800 6 io_oeb[1]
port 181 nsew signal output
rlabel metal2 s 181902 0 181958 800 6 io_oeb[20]
port 182 nsew signal output
rlabel metal2 s 189906 0 189962 800 6 io_oeb[21]
port 183 nsew signal output
rlabel metal2 s 197910 0 197966 800 6 io_oeb[22]
port 184 nsew signal output
rlabel metal2 s 205914 0 205970 800 6 io_oeb[23]
port 185 nsew signal output
rlabel metal2 s 213918 0 213974 800 6 io_oeb[24]
port 186 nsew signal output
rlabel metal2 s 221922 0 221978 800 6 io_oeb[25]
port 187 nsew signal output
rlabel metal2 s 229926 0 229982 800 6 io_oeb[26]
port 188 nsew signal output
rlabel metal2 s 237930 0 237986 800 6 io_oeb[27]
port 189 nsew signal output
rlabel metal2 s 245934 0 245990 800 6 io_oeb[28]
port 190 nsew signal output
rlabel metal2 s 253938 0 253994 800 6 io_oeb[29]
port 191 nsew signal output
rlabel metal2 s 37922 0 37978 800 6 io_oeb[2]
port 192 nsew signal output
rlabel metal2 s 261942 0 261998 800 6 io_oeb[30]
port 193 nsew signal output
rlabel metal2 s 269946 0 270002 800 6 io_oeb[31]
port 194 nsew signal output
rlabel metal2 s 277950 0 278006 800 6 io_oeb[32]
port 195 nsew signal output
rlabel metal2 s 281906 0 281962 800 6 io_oeb[33]
port 196 nsew signal output
rlabel metal2 s 285954 0 286010 800 6 io_oeb[34]
port 197 nsew signal output
rlabel metal2 s 289910 0 289966 800 6 io_oeb[35]
port 198 nsew signal output
rlabel metal2 s 293958 0 294014 800 6 io_oeb[36]
port 199 nsew signal output
rlabel metal2 s 297914 0 297970 800 6 io_oeb[37]
port 200 nsew signal output
rlabel metal2 s 45926 0 45982 800 6 io_oeb[3]
port 201 nsew signal output
rlabel metal2 s 53930 0 53986 800 6 io_oeb[4]
port 202 nsew signal output
rlabel metal2 s 61934 0 61990 800 6 io_oeb[5]
port 203 nsew signal output
rlabel metal2 s 69938 0 69994 800 6 io_oeb[6]
port 204 nsew signal output
rlabel metal2 s 77942 0 77998 800 6 io_oeb[7]
port 205 nsew signal output
rlabel metal2 s 85946 0 86002 800 6 io_oeb[8]
port 206 nsew signal output
rlabel metal2 s 93950 0 94006 800 6 io_oeb[9]
port 207 nsew signal output
rlabel metal2 s 25870 0 25926 800 6 io_ps[0]
port 208 nsew signal output
rlabel metal2 s 105910 0 105966 800 6 io_ps[10]
port 209 nsew signal output
rlabel metal2 s 113914 0 113970 800 6 io_ps[11]
port 210 nsew signal output
rlabel metal2 s 121918 0 121974 800 6 io_ps[12]
port 211 nsew signal output
rlabel metal2 s 129922 0 129978 800 6 io_ps[13]
port 212 nsew signal output
rlabel metal2 s 137926 0 137982 800 6 io_ps[14]
port 213 nsew signal output
rlabel metal2 s 145930 0 145986 800 6 io_ps[15]
port 214 nsew signal output
rlabel metal2 s 153934 0 153990 800 6 io_ps[16]
port 215 nsew signal output
rlabel metal2 s 161938 0 161994 800 6 io_ps[17]
port 216 nsew signal output
rlabel metal2 s 169942 0 169998 800 6 io_ps[18]
port 217 nsew signal output
rlabel metal2 s 177946 0 178002 800 6 io_ps[19]
port 218 nsew signal output
rlabel metal2 s 33874 0 33930 800 6 io_ps[1]
port 219 nsew signal output
rlabel metal2 s 185950 0 186006 800 6 io_ps[20]
port 220 nsew signal output
rlabel metal2 s 193954 0 194010 800 6 io_ps[21]
port 221 nsew signal output
rlabel metal2 s 201958 0 202014 800 6 io_ps[22]
port 222 nsew signal output
rlabel metal2 s 209870 0 209926 800 6 io_ps[23]
port 223 nsew signal output
rlabel metal2 s 217874 0 217930 800 6 io_ps[24]
port 224 nsew signal output
rlabel metal2 s 225878 0 225934 800 6 io_ps[25]
port 225 nsew signal output
rlabel metal2 s 233882 0 233938 800 6 io_ps[26]
port 226 nsew signal output
rlabel metal2 s 241886 0 241942 800 6 io_ps[27]
port 227 nsew signal output
rlabel metal2 s 249890 0 249946 800 6 io_ps[28]
port 228 nsew signal output
rlabel metal2 s 257894 0 257950 800 6 io_ps[29]
port 229 nsew signal output
rlabel metal2 s 41878 0 41934 800 6 io_ps[2]
port 230 nsew signal output
rlabel metal2 s 265898 0 265954 800 6 io_ps[30]
port 231 nsew signal output
rlabel metal2 s 273902 0 273958 800 6 io_ps[31]
port 232 nsew signal output
rlabel metal2 s 49882 0 49938 800 6 io_ps[3]
port 233 nsew signal output
rlabel metal2 s 57886 0 57942 800 6 io_ps[4]
port 234 nsew signal output
rlabel metal2 s 65890 0 65946 800 6 io_ps[5]
port 235 nsew signal output
rlabel metal2 s 73894 0 73950 800 6 io_ps[6]
port 236 nsew signal output
rlabel metal2 s 81898 0 81954 800 6 io_ps[7]
port 237 nsew signal output
rlabel metal2 s 89902 0 89958 800 6 io_ps[8]
port 238 nsew signal output
rlabel metal2 s 97906 0 97962 800 6 io_ps[9]
port 239 nsew signal output
rlabel metal2 s 5906 0 5962 800 6 rst_g
port 240 nsew signal input
rlabel metal2 s 13910 0 13966 800 6 rx
port 241 nsew signal input
rlabel metal2 s 9862 0 9918 800 6 tx
port 242 nsew signal output
rlabel metal3 s 0 3408 800 3528 6 vb_addr0[0]
port 243 nsew signal output
rlabel metal3 s 0 58080 800 58200 6 vb_addr0[10]
port 244 nsew signal output
rlabel metal3 s 0 63248 800 63368 6 vb_addr0[11]
port 245 nsew signal output
rlabel metal3 s 0 68280 800 68400 6 vb_addr0[12]
port 246 nsew signal output
rlabel metal3 s 0 9528 800 9648 6 vb_addr0[1]
port 247 nsew signal output
rlabel metal3 s 0 15512 800 15632 6 vb_addr0[2]
port 248 nsew signal output
rlabel metal3 s 0 21632 800 21752 6 vb_addr0[3]
port 249 nsew signal output
rlabel metal3 s 0 27752 800 27872 6 vb_addr0[4]
port 250 nsew signal output
rlabel metal3 s 0 32784 800 32904 6 vb_addr0[5]
port 251 nsew signal output
rlabel metal3 s 0 37816 800 37936 6 vb_addr0[6]
port 252 nsew signal output
rlabel metal3 s 0 42984 800 43104 6 vb_addr0[7]
port 253 nsew signal output
rlabel metal3 s 0 48016 800 48136 6 vb_addr0[8]
port 254 nsew signal output
rlabel metal3 s 0 53048 800 53168 6 vb_addr0[9]
port 255 nsew signal output
rlabel metal3 s 0 4360 800 4480 6 vb_addr1[0]
port 256 nsew signal output
rlabel metal3 s 0 59168 800 59288 6 vb_addr1[10]
port 257 nsew signal output
rlabel metal3 s 0 64200 800 64320 6 vb_addr1[11]
port 258 nsew signal output
rlabel metal3 s 0 69232 800 69352 6 vb_addr1[12]
port 259 nsew signal output
rlabel metal3 s 0 10480 800 10600 6 vb_addr1[1]
port 260 nsew signal output
rlabel metal3 s 0 16600 800 16720 6 vb_addr1[2]
port 261 nsew signal output
rlabel metal3 s 0 22584 800 22704 6 vb_addr1[3]
port 262 nsew signal output
rlabel metal3 s 0 28704 800 28824 6 vb_addr1[4]
port 263 nsew signal output
rlabel metal3 s 0 33736 800 33856 6 vb_addr1[5]
port 264 nsew signal output
rlabel metal3 s 0 38904 800 39024 6 vb_addr1[6]
port 265 nsew signal output
rlabel metal3 s 0 43936 800 44056 6 vb_addr1[7]
port 266 nsew signal output
rlabel metal3 s 0 48968 800 49088 6 vb_addr1[8]
port 267 nsew signal output
rlabel metal3 s 0 54000 800 54120 6 vb_addr1[9]
port 268 nsew signal output
rlabel metal3 s 0 416 800 536 6 vb_csb0
port 269 nsew signal output
rlabel metal3 s 0 1368 800 1488 6 vb_csb1
port 270 nsew signal output
rlabel metal3 s 0 5448 800 5568 6 vb_din0[0]
port 271 nsew signal output
rlabel metal3 s 0 60120 800 60240 6 vb_din0[10]
port 272 nsew signal output
rlabel metal3 s 0 65152 800 65272 6 vb_din0[11]
port 273 nsew signal output
rlabel metal3 s 0 70320 800 70440 6 vb_din0[12]
port 274 nsew signal output
rlabel metal3 s 0 73312 800 73432 6 vb_din0[13]
port 275 nsew signal output
rlabel metal3 s 0 76304 800 76424 6 vb_din0[14]
port 276 nsew signal output
rlabel metal3 s 0 79432 800 79552 6 vb_din0[15]
port 277 nsew signal output
rlabel metal3 s 0 82424 800 82544 6 vb_din0[16]
port 278 nsew signal output
rlabel metal3 s 0 85552 800 85672 6 vb_din0[17]
port 279 nsew signal output
rlabel metal3 s 0 88544 800 88664 6 vb_din0[18]
port 280 nsew signal output
rlabel metal3 s 0 91536 800 91656 6 vb_din0[19]
port 281 nsew signal output
rlabel metal3 s 0 11432 800 11552 6 vb_din0[1]
port 282 nsew signal output
rlabel metal3 s 0 94664 800 94784 6 vb_din0[20]
port 283 nsew signal output
rlabel metal3 s 0 97656 800 97776 6 vb_din0[21]
port 284 nsew signal output
rlabel metal3 s 0 100648 800 100768 6 vb_din0[22]
port 285 nsew signal output
rlabel metal3 s 0 103776 800 103896 6 vb_din0[23]
port 286 nsew signal output
rlabel metal3 s 0 106768 800 106888 6 vb_din0[24]
port 287 nsew signal output
rlabel metal3 s 0 109760 800 109880 6 vb_din0[25]
port 288 nsew signal output
rlabel metal3 s 0 112888 800 113008 6 vb_din0[26]
port 289 nsew signal output
rlabel metal3 s 0 115880 800 116000 6 vb_din0[27]
port 290 nsew signal output
rlabel metal3 s 0 118872 800 118992 6 vb_din0[28]
port 291 nsew signal output
rlabel metal3 s 0 122000 800 122120 6 vb_din0[29]
port 292 nsew signal output
rlabel metal3 s 0 17552 800 17672 6 vb_din0[2]
port 293 nsew signal output
rlabel metal3 s 0 124992 800 125112 6 vb_din0[30]
port 294 nsew signal output
rlabel metal3 s 0 128120 800 128240 6 vb_din0[31]
port 295 nsew signal output
rlabel metal3 s 0 23672 800 23792 6 vb_din0[3]
port 296 nsew signal output
rlabel metal3 s 0 29792 800 29912 6 vb_din0[4]
port 297 nsew signal output
rlabel metal3 s 0 34824 800 34944 6 vb_din0[5]
port 298 nsew signal output
rlabel metal3 s 0 39856 800 39976 6 vb_din0[6]
port 299 nsew signal output
rlabel metal3 s 0 44888 800 45008 6 vb_din0[7]
port 300 nsew signal output
rlabel metal3 s 0 50056 800 50176 6 vb_din0[8]
port 301 nsew signal output
rlabel metal3 s 0 55088 800 55208 6 vb_din0[9]
port 302 nsew signal output
rlabel metal3 s 0 6400 800 6520 6 vb_dout0[0]
port 303 nsew signal input
rlabel metal3 s 0 61208 800 61328 6 vb_dout0[10]
port 304 nsew signal input
rlabel metal3 s 0 66240 800 66360 6 vb_dout0[11]
port 305 nsew signal input
rlabel metal3 s 0 71272 800 71392 6 vb_dout0[12]
port 306 nsew signal input
rlabel metal3 s 0 74400 800 74520 6 vb_dout0[13]
port 307 nsew signal input
rlabel metal3 s 0 77392 800 77512 6 vb_dout0[14]
port 308 nsew signal input
rlabel metal3 s 0 80384 800 80504 6 vb_dout0[15]
port 309 nsew signal input
rlabel metal3 s 0 83512 800 83632 6 vb_dout0[16]
port 310 nsew signal input
rlabel metal3 s 0 86504 800 86624 6 vb_dout0[17]
port 311 nsew signal input
rlabel metal3 s 0 89496 800 89616 6 vb_dout0[18]
port 312 nsew signal input
rlabel metal3 s 0 92624 800 92744 6 vb_dout0[19]
port 313 nsew signal input
rlabel metal3 s 0 12520 800 12640 6 vb_dout0[1]
port 314 nsew signal input
rlabel metal3 s 0 95616 800 95736 6 vb_dout0[20]
port 315 nsew signal input
rlabel metal3 s 0 98608 800 98728 6 vb_dout0[21]
port 316 nsew signal input
rlabel metal3 s 0 101736 800 101856 6 vb_dout0[22]
port 317 nsew signal input
rlabel metal3 s 0 104728 800 104848 6 vb_dout0[23]
port 318 nsew signal input
rlabel metal3 s 0 107720 800 107840 6 vb_dout0[24]
port 319 nsew signal input
rlabel metal3 s 0 110848 800 110968 6 vb_dout0[25]
port 320 nsew signal input
rlabel metal3 s 0 113840 800 113960 6 vb_dout0[26]
port 321 nsew signal input
rlabel metal3 s 0 116968 800 117088 6 vb_dout0[27]
port 322 nsew signal input
rlabel metal3 s 0 119960 800 120080 6 vb_dout0[28]
port 323 nsew signal input
rlabel metal3 s 0 122952 800 123072 6 vb_dout0[29]
port 324 nsew signal input
rlabel metal3 s 0 18640 800 18760 6 vb_dout0[2]
port 325 nsew signal input
rlabel metal3 s 0 126080 800 126200 6 vb_dout0[30]
port 326 nsew signal input
rlabel metal3 s 0 129072 800 129192 6 vb_dout0[31]
port 327 nsew signal input
rlabel metal3 s 0 24624 800 24744 6 vb_dout0[3]
port 328 nsew signal input
rlabel metal3 s 0 30744 800 30864 6 vb_dout0[4]
port 329 nsew signal input
rlabel metal3 s 0 35776 800 35896 6 vb_dout0[5]
port 330 nsew signal input
rlabel metal3 s 0 40944 800 41064 6 vb_dout0[6]
port 331 nsew signal input
rlabel metal3 s 0 45976 800 46096 6 vb_dout0[7]
port 332 nsew signal input
rlabel metal3 s 0 51008 800 51128 6 vb_dout0[8]
port 333 nsew signal input
rlabel metal3 s 0 56040 800 56160 6 vb_dout0[9]
port 334 nsew signal input
rlabel metal3 s 0 7488 800 7608 6 vb_dout1[0]
port 335 nsew signal input
rlabel metal3 s 0 62160 800 62280 6 vb_dout1[10]
port 336 nsew signal input
rlabel metal3 s 0 67192 800 67312 6 vb_dout1[11]
port 337 nsew signal input
rlabel metal3 s 0 72360 800 72480 6 vb_dout1[12]
port 338 nsew signal input
rlabel metal3 s 0 75352 800 75472 6 vb_dout1[13]
port 339 nsew signal input
rlabel metal3 s 0 78344 800 78464 6 vb_dout1[14]
port 340 nsew signal input
rlabel metal3 s 0 81472 800 81592 6 vb_dout1[15]
port 341 nsew signal input
rlabel metal3 s 0 84464 800 84584 6 vb_dout1[16]
port 342 nsew signal input
rlabel metal3 s 0 87456 800 87576 6 vb_dout1[17]
port 343 nsew signal input
rlabel metal3 s 0 90584 800 90704 6 vb_dout1[18]
port 344 nsew signal input
rlabel metal3 s 0 93576 800 93696 6 vb_dout1[19]
port 345 nsew signal input
rlabel metal3 s 0 13472 800 13592 6 vb_dout1[1]
port 346 nsew signal input
rlabel metal3 s 0 96704 800 96824 6 vb_dout1[20]
port 347 nsew signal input
rlabel metal3 s 0 99696 800 99816 6 vb_dout1[21]
port 348 nsew signal input
rlabel metal3 s 0 102688 800 102808 6 vb_dout1[22]
port 349 nsew signal input
rlabel metal3 s 0 105816 800 105936 6 vb_dout1[23]
port 350 nsew signal input
rlabel metal3 s 0 108808 800 108928 6 vb_dout1[24]
port 351 nsew signal input
rlabel metal3 s 0 111800 800 111920 6 vb_dout1[25]
port 352 nsew signal input
rlabel metal3 s 0 114928 800 115048 6 vb_dout1[26]
port 353 nsew signal input
rlabel metal3 s 0 117920 800 118040 6 vb_dout1[27]
port 354 nsew signal input
rlabel metal3 s 0 120912 800 121032 6 vb_dout1[28]
port 355 nsew signal input
rlabel metal3 s 0 124040 800 124160 6 vb_dout1[29]
port 356 nsew signal input
rlabel metal3 s 0 19592 800 19712 6 vb_dout1[2]
port 357 nsew signal input
rlabel metal3 s 0 127032 800 127152 6 vb_dout1[30]
port 358 nsew signal input
rlabel metal3 s 0 130024 800 130144 6 vb_dout1[31]
port 359 nsew signal input
rlabel metal3 s 0 25712 800 25832 6 vb_dout1[3]
port 360 nsew signal input
rlabel metal3 s 0 31832 800 31952 6 vb_dout1[4]
port 361 nsew signal input
rlabel metal3 s 0 36864 800 36984 6 vb_dout1[5]
port 362 nsew signal input
rlabel metal3 s 0 41896 800 42016 6 vb_dout1[6]
port 363 nsew signal input
rlabel metal3 s 0 46928 800 47048 6 vb_dout1[7]
port 364 nsew signal input
rlabel metal3 s 0 52096 800 52216 6 vb_dout1[8]
port 365 nsew signal input
rlabel metal3 s 0 57128 800 57248 6 vb_dout1[9]
port 366 nsew signal input
rlabel metal3 s 0 2320 800 2440 6 vb_web0
port 367 nsew signal output
rlabel metal3 s 0 8440 800 8560 6 vb_wmask0[0]
port 368 nsew signal output
rlabel metal3 s 0 14560 800 14680 6 vb_wmask0[1]
port 369 nsew signal output
rlabel metal3 s 0 20680 800 20800 6 vb_wmask0[2]
port 370 nsew signal output
rlabel metal3 s 0 26664 800 26784 6 vb_wmask0[3]
port 371 nsew signal output
rlabel metal4 s 4208 2128 4528 297616 6 vccd1
port 372 nsew power input
rlabel metal4 s 34928 2128 35248 297616 6 vccd1
port 372 nsew power input
rlabel metal4 s 65648 2128 65968 297616 6 vccd1
port 372 nsew power input
rlabel metal4 s 96368 2128 96688 297616 6 vccd1
port 372 nsew power input
rlabel metal4 s 127088 2128 127408 297616 6 vccd1
port 372 nsew power input
rlabel metal4 s 157808 2128 158128 297616 6 vccd1
port 372 nsew power input
rlabel metal4 s 188528 2128 188848 297616 6 vccd1
port 372 nsew power input
rlabel metal4 s 219248 2128 219568 297616 6 vccd1
port 372 nsew power input
rlabel metal4 s 249968 2128 250288 297616 6 vccd1
port 372 nsew power input
rlabel metal4 s 280688 2128 281008 297616 6 vccd1
port 372 nsew power input
rlabel metal4 s 19568 2128 19888 297616 6 vssd1
port 373 nsew ground input
rlabel metal4 s 50288 2128 50608 297616 6 vssd1
port 373 nsew ground input
rlabel metal4 s 81008 2128 81328 297616 6 vssd1
port 373 nsew ground input
rlabel metal4 s 111728 2128 112048 297616 6 vssd1
port 373 nsew ground input
rlabel metal4 s 142448 2128 142768 297616 6 vssd1
port 373 nsew ground input
rlabel metal4 s 173168 2128 173488 297616 6 vssd1
port 373 nsew ground input
rlabel metal4 s 203888 2128 204208 297616 6 vssd1
port 373 nsew ground input
rlabel metal4 s 234608 2128 234928 297616 6 vssd1
port 373 nsew ground input
rlabel metal4 s 265328 2128 265648 297616 6 vssd1
port 373 nsew ground input
rlabel metal4 s 296048 2128 296368 297616 6 vssd1
port 373 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 300000 300000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 76529094
string GDS_FILE /home/kasirga/c0_hayyan/GL_GECTI/caravel_user_project/openlane/c0_system/runs/c0_system/results/finishing/c0_system.magic.gds
string GDS_START 1666336
<< end >>


magic
tech sky130A
magscale 1 2
timestamp 1647512816
<< metal1 >>
rect 154114 700476 154120 700528
rect 154172 700516 154178 700528
rect 233878 700516 233884 700528
rect 154172 700488 233884 700516
rect 154172 700476 154178 700488
rect 233878 700476 233884 700488
rect 233936 700476 233942 700528
rect 89162 700408 89168 700460
rect 89220 700448 89226 700460
rect 191098 700448 191104 700460
rect 89220 700420 191104 700448
rect 89220 700408 89226 700420
rect 191098 700408 191104 700420
rect 191156 700408 191162 700460
rect 202782 700408 202788 700460
rect 202840 700448 202846 700460
rect 239398 700448 239404 700460
rect 202840 700420 239404 700448
rect 202840 700408 202846 700420
rect 239398 700408 239404 700420
rect 239456 700408 239462 700460
rect 137830 700340 137836 700392
rect 137888 700380 137894 700392
rect 239582 700380 239588 700392
rect 137888 700352 239588 700380
rect 137888 700340 137894 700352
rect 239582 700340 239588 700352
rect 239640 700340 239646 700392
rect 262214 700340 262220 700392
rect 262272 700380 262278 700392
rect 332502 700380 332508 700392
rect 262272 700352 332508 700380
rect 262272 700340 262278 700352
rect 332502 700340 332508 700352
rect 332560 700340 332566 700392
rect 72970 700272 72976 700324
rect 73028 700312 73034 700324
rect 239490 700312 239496 700324
rect 73028 700284 239496 700312
rect 73028 700272 73034 700284
rect 239490 700272 239496 700284
rect 239548 700272 239554 700324
rect 262122 700272 262128 700324
rect 262180 700312 262186 700324
rect 348786 700312 348792 700324
rect 262180 700284 348792 700312
rect 262180 700272 262186 700284
rect 348786 700272 348792 700284
rect 348844 700272 348850 700324
rect 500218 700272 500224 700324
rect 500276 700312 500282 700324
rect 527174 700312 527180 700324
rect 500276 700284 527180 700312
rect 500276 700272 500282 700284
rect 527174 700272 527180 700284
rect 527232 700272 527238 700324
rect 397454 699660 397460 699712
rect 397512 699700 397518 699712
rect 403618 699700 403624 699712
rect 397512 699672 403624 699700
rect 397512 699660 397518 699672
rect 403618 699660 403624 699672
rect 403676 699660 403682 699712
rect 413646 698096 413652 698148
rect 413704 698136 413710 698148
rect 416038 698136 416044 698148
rect 413704 698108 416044 698136
rect 413704 698096 413710 698108
rect 416038 698096 416044 698108
rect 416096 698096 416102 698148
rect 266354 697552 266360 697604
rect 266412 697592 266418 697604
rect 267642 697592 267648 697604
rect 266412 697564 267648 697592
rect 266412 697552 266418 697564
rect 267642 697552 267648 697564
rect 267700 697552 267706 697604
rect 261938 696940 261944 696992
rect 261996 696980 262002 696992
rect 262214 696980 262220 696992
rect 261996 696952 262220 696980
rect 261996 696940 262002 696952
rect 262214 696940 262220 696952
rect 262272 696940 262278 696992
rect 259454 694084 259460 694136
rect 259512 694124 259518 694136
rect 261938 694124 261944 694136
rect 259512 694096 261944 694124
rect 259512 694084 259518 694096
rect 261938 694084 261944 694096
rect 261996 694084 262002 694136
rect 259546 694016 259552 694068
rect 259604 694056 259610 694068
rect 262122 694056 262128 694068
rect 259604 694028 262128 694056
rect 259604 694016 259610 694028
rect 262122 694016 262128 694028
rect 262180 694016 262186 694068
rect 257338 691364 257344 691416
rect 257396 691404 257402 691416
rect 259546 691404 259552 691416
rect 257396 691376 259552 691404
rect 257396 691364 257402 691376
rect 259546 691364 259552 691376
rect 259604 691364 259610 691416
rect 403618 687148 403624 687200
rect 403676 687188 403682 687200
rect 406378 687188 406384 687200
rect 403676 687160 406384 687188
rect 403676 687148 403682 687160
rect 406378 687148 406384 687160
rect 406436 687148 406442 687200
rect 253198 683136 253204 683188
rect 253256 683176 253262 683188
rect 259362 683176 259368 683188
rect 253256 683148 259368 683176
rect 253256 683136 253262 683148
rect 259362 683136 259368 683148
rect 259420 683136 259426 683188
rect 3418 671032 3424 671084
rect 3476 671072 3482 671084
rect 7558 671072 7564 671084
rect 3476 671044 7564 671072
rect 3476 671032 3482 671044
rect 7558 671032 7564 671044
rect 7616 671032 7622 671084
rect 256050 668584 256056 668636
rect 256108 668624 256114 668636
rect 257338 668624 257344 668636
rect 256108 668596 257344 668624
rect 256108 668584 256114 668596
rect 257338 668584 257344 668596
rect 257396 668584 257402 668636
rect 254578 664912 254584 664964
rect 254636 664952 254642 664964
rect 256050 664952 256056 664964
rect 254636 664924 256056 664952
rect 254636 664912 254642 664924
rect 256050 664912 256056 664924
rect 256108 664912 256114 664964
rect 3418 656888 3424 656940
rect 3476 656928 3482 656940
rect 233970 656928 233976 656940
rect 3476 656900 233976 656928
rect 3476 656888 3482 656900
rect 233970 656888 233976 656900
rect 234028 656888 234034 656940
rect 416038 655460 416044 655512
rect 416096 655500 416102 655512
rect 419442 655500 419448 655512
rect 416096 655472 419448 655500
rect 416096 655460 416102 655472
rect 419442 655460 419448 655472
rect 419500 655460 419506 655512
rect 419442 651312 419448 651364
rect 419500 651352 419506 651364
rect 424318 651352 424324 651364
rect 419500 651324 424324 651352
rect 419500 651312 419506 651324
rect 424318 651312 424324 651324
rect 424376 651312 424382 651364
rect 406378 647164 406384 647216
rect 406436 647204 406442 647216
rect 409138 647204 409144 647216
rect 406436 647176 409144 647204
rect 406436 647164 406442 647176
rect 409138 647164 409144 647176
rect 409196 647164 409202 647216
rect 424318 638188 424324 638240
rect 424376 638228 424382 638240
rect 432598 638228 432604 638240
rect 424376 638200 432604 638228
rect 424376 638188 424382 638200
rect 432598 638188 432604 638200
rect 432656 638188 432662 638240
rect 409138 636828 409144 636880
rect 409196 636868 409202 636880
rect 414014 636868 414020 636880
rect 409196 636840 414020 636868
rect 409196 636828 409202 636840
rect 414014 636828 414020 636840
rect 414072 636828 414078 636880
rect 414014 634040 414020 634092
rect 414072 634080 414078 634092
rect 424134 634080 424140 634092
rect 414072 634052 424140 634080
rect 414072 634040 414078 634052
rect 424134 634040 424140 634052
rect 424192 634040 424198 634092
rect 424134 628532 424140 628584
rect 424192 628572 424198 628584
rect 447778 628572 447784 628584
rect 424192 628544 447784 628572
rect 424192 628532 424198 628544
rect 447778 628532 447784 628544
rect 447836 628532 447842 628584
rect 253290 619556 253296 619608
rect 253348 619596 253354 619608
rect 254578 619596 254584 619608
rect 253348 619568 254584 619596
rect 253348 619556 253354 619568
rect 254578 619556 254584 619568
rect 254636 619556 254642 619608
rect 251818 610444 251824 610496
rect 251876 610484 251882 610496
rect 253290 610484 253296 610496
rect 251876 610456 253296 610484
rect 251876 610444 251882 610456
rect 253290 610444 253296 610456
rect 253348 610444 253354 610496
rect 432598 609220 432604 609272
rect 432656 609260 432662 609272
rect 442258 609260 442264 609272
rect 432656 609232 442264 609260
rect 432656 609220 432662 609232
rect 442258 609220 442264 609232
rect 442316 609220 442322 609272
rect 3510 605820 3516 605872
rect 3568 605860 3574 605872
rect 239674 605860 239680 605872
rect 3568 605832 239680 605860
rect 3568 605820 3574 605832
rect 239674 605820 239680 605832
rect 239732 605820 239738 605872
rect 447778 591948 447784 592000
rect 447836 591988 447842 592000
rect 453298 591988 453304 592000
rect 447836 591960 453304 591988
rect 447836 591948 447842 591960
rect 453298 591948 453304 591960
rect 453356 591948 453362 592000
rect 251818 590696 251824 590708
rect 249812 590668 251824 590696
rect 249058 590588 249064 590640
rect 249116 590628 249122 590640
rect 249812 590628 249840 590668
rect 251818 590656 251824 590668
rect 251876 590656 251882 590708
rect 249116 590600 249840 590628
rect 249116 590588 249122 590600
rect 442258 579572 442264 579624
rect 442316 579612 442322 579624
rect 445662 579612 445668 579624
rect 442316 579584 445668 579612
rect 442316 579572 442322 579584
rect 445662 579572 445668 579584
rect 445720 579572 445726 579624
rect 445662 574200 445668 574252
rect 445720 574240 445726 574252
rect 447778 574240 447784 574252
rect 445720 574212 447784 574240
rect 445720 574200 445726 574212
rect 447778 574200 447784 574212
rect 447836 574200 447842 574252
rect 251818 563048 251824 563100
rect 251876 563088 251882 563100
rect 253198 563088 253204 563100
rect 251876 563060 253204 563088
rect 251876 563048 251882 563060
rect 253198 563048 253204 563060
rect 253256 563048 253262 563100
rect 453298 562300 453304 562352
rect 453356 562340 453362 562352
rect 456058 562340 456064 562352
rect 453356 562312 456064 562340
rect 453356 562300 453362 562312
rect 456058 562300 456064 562312
rect 456116 562300 456122 562352
rect 447778 559716 447784 559768
rect 447836 559756 447842 559768
rect 451274 559756 451280 559768
rect 447836 559728 451280 559756
rect 447836 559716 447842 559728
rect 451274 559716 451280 559728
rect 451332 559716 451338 559768
rect 451274 556792 451280 556844
rect 451332 556832 451338 556844
rect 461670 556832 461676 556844
rect 451332 556804 461676 556832
rect 451332 556792 451338 556804
rect 461670 556792 461676 556804
rect 461728 556792 461734 556844
rect 456058 554684 456064 554736
rect 456116 554724 456122 554736
rect 461578 554724 461584 554736
rect 456116 554696 461584 554724
rect 456116 554684 456122 554696
rect 461578 554684 461584 554696
rect 461636 554684 461642 554736
rect 461670 554684 461676 554736
rect 461728 554724 461734 554736
rect 465718 554724 465724 554736
rect 461728 554696 465724 554724
rect 461728 554684 461734 554696
rect 465718 554684 465724 554696
rect 465776 554684 465782 554736
rect 3602 553392 3608 553444
rect 3660 553432 3666 553444
rect 239766 553432 239772 553444
rect 3660 553404 239772 553432
rect 3660 553392 3666 553404
rect 239766 553392 239772 553404
rect 239824 553392 239830 553444
rect 260098 540200 260104 540252
rect 260156 540240 260162 540252
rect 282914 540240 282920 540252
rect 260156 540212 282920 540240
rect 260156 540200 260162 540212
rect 282914 540200 282920 540212
rect 282972 540200 282978 540252
rect 461578 538840 461584 538892
rect 461636 538880 461642 538892
rect 472618 538880 472624 538892
rect 461636 538852 472624 538880
rect 461636 538840 461642 538852
rect 472618 538840 472624 538852
rect 472676 538840 472682 538892
rect 465718 534692 465724 534744
rect 465776 534732 465782 534744
rect 475470 534732 475476 534744
rect 465776 534704 475476 534732
rect 465776 534692 465782 534704
rect 475470 534692 475476 534704
rect 475528 534692 475534 534744
rect 472618 529864 472624 529916
rect 472676 529904 472682 529916
rect 475378 529904 475384 529916
rect 472676 529876 475384 529904
rect 472676 529864 472682 529876
rect 475378 529864 475384 529876
rect 475436 529864 475442 529916
rect 475470 526668 475476 526720
rect 475528 526708 475534 526720
rect 479518 526708 479524 526720
rect 475528 526680 479524 526708
rect 475528 526668 475534 526680
rect 479518 526668 479524 526680
rect 479576 526668 479582 526720
rect 258718 525784 258724 525836
rect 258776 525824 258782 525836
rect 260098 525824 260104 525836
rect 258776 525796 260104 525824
rect 258776 525784 258782 525796
rect 260098 525784 260104 525796
rect 260156 525784 260162 525836
rect 249426 524424 249432 524476
rect 249484 524464 249490 524476
rect 251818 524464 251824 524476
rect 249484 524436 251824 524464
rect 249484 524424 249490 524436
rect 251818 524424 251824 524436
rect 251876 524424 251882 524476
rect 498838 524424 498844 524476
rect 498896 524464 498902 524476
rect 580166 524464 580172 524476
rect 498896 524436 580172 524464
rect 498896 524424 498902 524436
rect 580166 524424 580172 524436
rect 580224 524424 580230 524476
rect 247678 520276 247684 520328
rect 247736 520316 247742 520328
rect 249426 520316 249432 520328
rect 247736 520288 249432 520316
rect 247736 520276 247742 520288
rect 249426 520276 249432 520288
rect 249484 520276 249490 520328
rect 479518 514020 479524 514072
rect 479576 514060 479582 514072
rect 490558 514060 490564 514072
rect 479576 514032 490564 514060
rect 479576 514020 479582 514032
rect 490558 514020 490564 514032
rect 490616 514020 490622 514072
rect 257338 506676 257344 506728
rect 257396 506716 257402 506728
rect 258718 506716 258724 506728
rect 257396 506688 258724 506716
rect 257396 506676 257402 506688
rect 258718 506676 258724 506688
rect 258776 506676 258782 506728
rect 246298 503616 246304 503668
rect 246356 503656 246362 503668
rect 249058 503656 249064 503668
rect 246356 503628 249064 503656
rect 246356 503616 246362 503628
rect 249058 503616 249064 503628
rect 249116 503616 249122 503668
rect 2866 500964 2872 501016
rect 2924 501004 2930 501016
rect 239858 501004 239864 501016
rect 2924 500976 239864 501004
rect 2924 500964 2930 500976
rect 239858 500964 239864 500976
rect 239916 500964 239922 501016
rect 253934 496816 253940 496868
rect 253992 496856 253998 496868
rect 257338 496856 257344 496868
rect 253992 496828 257344 496856
rect 253992 496816 253998 496828
rect 257338 496816 257344 496828
rect 257396 496816 257402 496868
rect 247770 490560 247776 490612
rect 247828 490600 247834 490612
rect 253934 490600 253940 490612
rect 247828 490572 253940 490600
rect 247828 490560 247834 490572
rect 253934 490560 253940 490572
rect 253992 490560 253998 490612
rect 244918 473968 244924 474020
rect 244976 474008 244982 474020
rect 247770 474008 247776 474020
rect 244976 473980 247776 474008
rect 244976 473968 244982 473980
rect 247770 473968 247776 473980
rect 247828 473968 247834 474020
rect 113818 466012 113824 466064
rect 113876 466052 113882 466064
rect 238018 466052 238024 466064
rect 113876 466024 238024 466052
rect 113876 466012 113882 466024
rect 238018 466012 238024 466024
rect 238076 466012 238082 466064
rect 169754 465944 169760 465996
rect 169812 465984 169818 465996
rect 192478 465984 192484 465996
rect 169812 465956 192484 465984
rect 169812 465944 169818 465956
rect 192478 465944 192484 465956
rect 192536 465944 192542 465996
rect 156138 465876 156144 465928
rect 156196 465916 156202 465928
rect 186774 465916 186780 465928
rect 156196 465888 186780 465916
rect 156196 465876 156202 465888
rect 186774 465876 186780 465888
rect 186832 465876 186838 465928
rect 153378 465808 153384 465860
rect 153436 465848 153442 465860
rect 186682 465848 186688 465860
rect 153436 465820 186688 465848
rect 153436 465808 153442 465820
rect 186682 465808 186688 465820
rect 186740 465808 186746 465860
rect 136082 465740 136088 465792
rect 136140 465780 136146 465792
rect 192662 465780 192668 465792
rect 136140 465752 192668 465780
rect 136140 465740 136146 465752
rect 192662 465740 192668 465752
rect 192720 465740 192726 465792
rect 128722 465672 128728 465724
rect 128780 465712 128786 465724
rect 187142 465712 187148 465724
rect 128780 465684 187148 465712
rect 128780 465672 128786 465684
rect 187142 465672 187148 465684
rect 187200 465672 187206 465724
rect 91186 465604 91192 465656
rect 91244 465644 91250 465656
rect 168374 465644 168380 465656
rect 91244 465616 168380 465644
rect 91244 465604 91250 465616
rect 168374 465604 168380 465616
rect 168432 465604 168438 465656
rect 168466 465604 168472 465656
rect 168524 465644 168530 465656
rect 192570 465644 192576 465656
rect 168524 465616 192576 465644
rect 168524 465604 168530 465616
rect 192570 465604 192576 465616
rect 192628 465604 192634 465656
rect 111058 465536 111064 465588
rect 111116 465576 111122 465588
rect 188430 465576 188436 465588
rect 111116 465548 188436 465576
rect 111116 465536 111122 465548
rect 188430 465536 188436 465548
rect 188488 465536 188494 465588
rect 101674 465468 101680 465520
rect 101732 465508 101738 465520
rect 189718 465508 189724 465520
rect 101732 465480 189724 465508
rect 101732 465468 101738 465480
rect 189718 465468 189724 465480
rect 189776 465468 189782 465520
rect 103698 465400 103704 465452
rect 103756 465440 103762 465452
rect 193858 465440 193864 465452
rect 103756 465412 193864 465440
rect 103756 465400 103762 465412
rect 193858 465400 193864 465412
rect 193916 465400 193922 465452
rect 98546 465332 98552 465384
rect 98604 465372 98610 465384
rect 198090 465372 198096 465384
rect 98604 465344 198096 465372
rect 98604 465332 98610 465344
rect 198090 465332 198096 465344
rect 198148 465332 198154 465384
rect 96154 465264 96160 465316
rect 96212 465304 96218 465316
rect 197998 465304 198004 465316
rect 96212 465276 198004 465304
rect 96212 465264 96218 465276
rect 197998 465264 198004 465276
rect 198056 465264 198062 465316
rect 118602 465196 118608 465248
rect 118660 465236 118666 465248
rect 238202 465236 238208 465248
rect 118660 465208 238208 465236
rect 118660 465196 118666 465208
rect 238202 465196 238208 465208
rect 238260 465196 238266 465248
rect 116210 465128 116216 465180
rect 116268 465168 116274 465180
rect 238110 465168 238116 465180
rect 116268 465140 238116 465168
rect 116268 465128 116274 465140
rect 238110 465128 238116 465140
rect 238168 465128 238174 465180
rect 143626 465060 143632 465112
rect 143684 465100 143690 465112
rect 155862 465100 155868 465112
rect 143684 465072 155868 465100
rect 143684 465060 143690 465072
rect 155862 465060 155868 465072
rect 155920 465060 155926 465112
rect 141050 464992 141056 465044
rect 141108 465032 141114 465044
rect 191282 465032 191288 465044
rect 141108 465004 191288 465032
rect 141108 464992 141114 465004
rect 191282 464992 191288 465004
rect 191340 464992 191346 465044
rect 133506 464924 133512 464976
rect 133564 464964 133570 464976
rect 188706 464964 188712 464976
rect 133564 464936 188712 464964
rect 133564 464924 133570 464936
rect 188706 464924 188712 464936
rect 188764 464924 188770 464976
rect 179414 464856 179420 464908
rect 179472 464896 179478 464908
rect 235258 464896 235264 464908
rect 179472 464868 235264 464896
rect 179472 464856 179478 464868
rect 235258 464856 235264 464868
rect 235316 464856 235322 464908
rect 131114 464788 131120 464840
rect 131172 464828 131178 464840
rect 188614 464828 188620 464840
rect 131172 464800 188620 464828
rect 131172 464788 131178 464800
rect 188614 464788 188620 464800
rect 188672 464788 188678 464840
rect 125962 464720 125968 464772
rect 126020 464760 126026 464772
rect 188522 464760 188528 464772
rect 126020 464732 188528 464760
rect 126020 464720 126026 464732
rect 188522 464720 188528 464732
rect 188580 464720 188586 464772
rect 123570 464652 123576 464704
rect 123628 464692 123634 464704
rect 187050 464692 187056 464704
rect 123628 464664 187056 464692
rect 123628 464652 123634 464664
rect 187050 464652 187056 464664
rect 187108 464652 187114 464704
rect 120994 464584 121000 464636
rect 121052 464624 121058 464636
rect 186958 464624 186964 464636
rect 121052 464596 186964 464624
rect 121052 464584 121058 464596
rect 186958 464584 186964 464596
rect 187016 464584 187022 464636
rect 168374 464516 168380 464568
rect 168432 464556 168438 464568
rect 235350 464556 235356 464568
rect 168432 464528 235356 464556
rect 168432 464516 168438 464528
rect 235350 464516 235356 464528
rect 235408 464516 235414 464568
rect 155862 464448 155868 464500
rect 155920 464488 155926 464500
rect 238386 464488 238392 464500
rect 155920 464460 238392 464488
rect 155920 464448 155926 464460
rect 238386 464448 238392 464460
rect 238444 464448 238450 464500
rect 138474 464380 138480 464432
rect 138532 464420 138538 464432
rect 238294 464420 238300 464432
rect 138532 464392 238300 464420
rect 138532 464380 138538 464392
rect 238294 464380 238300 464392
rect 238352 464380 238358 464432
rect 83458 464312 83464 464364
rect 83516 464352 83522 464364
rect 196618 464352 196624 464364
rect 83516 464324 196624 464352
rect 83516 464312 83522 464324
rect 196618 464312 196624 464324
rect 196676 464312 196682 464364
rect 146018 464244 146024 464296
rect 146076 464284 146082 464296
rect 191466 464284 191472 464296
rect 146076 464256 191472 464284
rect 146076 464244 146082 464256
rect 191466 464244 191472 464256
rect 191524 464244 191530 464296
rect 148502 464176 148508 464228
rect 148560 464216 148566 464228
rect 191374 464216 191380 464228
rect 148560 464188 191380 464216
rect 148560 464176 148566 464188
rect 191374 464176 191380 464188
rect 191432 464176 191438 464228
rect 151078 464108 151084 464160
rect 151136 464148 151142 464160
rect 189902 464148 189908 464160
rect 151136 464120 189908 464148
rect 151136 464108 151142 464120
rect 189902 464108 189908 464120
rect 189960 464108 189966 464160
rect 186682 463020 186688 463072
rect 186740 463060 186746 463072
rect 238478 463060 238484 463072
rect 186740 463032 238484 463060
rect 186740 463020 186746 463032
rect 238478 463020 238484 463032
rect 238536 463020 238542 463072
rect 186774 462952 186780 463004
rect 186832 462992 186838 463004
rect 238570 462992 238576 463004
rect 186832 462964 238576 462992
rect 186832 462952 186838 462964
rect 238570 462952 238576 462964
rect 238628 462952 238634 463004
rect 189074 458192 189080 458244
rect 189132 458232 189138 458244
rect 195330 458232 195336 458244
rect 189132 458204 195336 458232
rect 189132 458192 189138 458204
rect 195330 458192 195336 458204
rect 195388 458192 195394 458244
rect 245010 455336 245016 455388
rect 245068 455376 245074 455388
rect 247678 455376 247684 455388
rect 245068 455348 247684 455376
rect 245068 455336 245074 455348
rect 247678 455336 247684 455348
rect 247736 455336 247742 455388
rect 245102 452548 245108 452600
rect 245160 452588 245166 452600
rect 246298 452588 246304 452600
rect 245160 452560 246304 452588
rect 245160 452548 245166 452560
rect 246298 452548 246304 452560
rect 246356 452548 246362 452600
rect 2958 448536 2964 448588
rect 3016 448576 3022 448588
rect 43438 448576 43444 448588
rect 3016 448548 43444 448576
rect 3016 448536 3022 448548
rect 43438 448536 43444 448548
rect 43496 448536 43502 448588
rect 242526 445816 242532 445868
rect 242584 445856 242590 445868
rect 245010 445856 245016 445868
rect 242584 445828 245016 445856
rect 242584 445816 242590 445828
rect 245010 445816 245016 445828
rect 245068 445816 245074 445868
rect 242894 444456 242900 444508
rect 242952 444496 242958 444508
rect 244918 444496 244924 444508
rect 242952 444468 244924 444496
rect 242952 444456 242958 444468
rect 244918 444456 244924 444468
rect 244976 444456 244982 444508
rect 240226 443368 240232 443420
rect 240284 443408 240290 443420
rect 245102 443408 245108 443420
rect 240284 443380 245108 443408
rect 240284 443368 240290 443380
rect 245102 443368 245108 443380
rect 245160 443368 245166 443420
rect 240134 442416 240140 442468
rect 240192 442456 240198 442468
rect 242526 442456 242532 442468
rect 240192 442428 242532 442456
rect 240192 442416 240198 442428
rect 242526 442416 242532 442428
rect 242584 442416 242590 442468
rect 242066 442280 242072 442332
rect 242124 442320 242130 442332
rect 242894 442320 242900 442332
rect 242124 442292 242900 442320
rect 242124 442280 242130 442292
rect 242894 442280 242900 442292
rect 242952 442280 242958 442332
rect 240042 440852 240048 440904
rect 240100 440892 240106 440904
rect 266354 440892 266360 440904
rect 240100 440864 266360 440892
rect 240100 440852 240106 440864
rect 266354 440852 266360 440864
rect 266412 440852 266418 440904
rect 240410 440240 240416 440292
rect 240468 440280 240474 440292
rect 242066 440280 242072 440292
rect 240468 440252 242072 440280
rect 240468 440240 240474 440252
rect 242066 440240 242072 440252
rect 242124 440240 242130 440292
rect 239950 438880 239956 438932
rect 240008 438920 240014 438932
rect 240134 438920 240140 438932
rect 240008 438892 240140 438920
rect 240008 438880 240014 438892
rect 240134 438880 240140 438892
rect 240192 438880 240198 438932
rect 198182 437520 198188 437572
rect 198240 437560 198246 437572
rect 237466 437560 237472 437572
rect 198240 437532 237472 437560
rect 198240 437520 198246 437532
rect 237466 437520 237472 437532
rect 237524 437520 237530 437572
rect 189810 437452 189816 437504
rect 189868 437492 189874 437504
rect 237374 437492 237380 437504
rect 189868 437464 237380 437492
rect 189868 437452 189874 437464
rect 237374 437452 237380 437464
rect 237432 437452 237438 437504
rect 239306 436568 239312 436620
rect 239364 436608 239370 436620
rect 240226 436608 240232 436620
rect 239364 436580 240232 436608
rect 239364 436568 239370 436580
rect 240226 436568 240232 436580
rect 240284 436568 240290 436620
rect 191190 433372 191196 433424
rect 191248 433412 191254 433424
rect 237374 433412 237380 433424
rect 191248 433384 237380 433412
rect 191248 433372 191254 433384
rect 237374 433372 237380 433384
rect 237432 433372 237438 433424
rect 188798 433304 188804 433356
rect 188856 433344 188862 433356
rect 237466 433344 237472 433356
rect 188856 433316 237472 433344
rect 188856 433304 188862 433316
rect 237466 433304 237472 433316
rect 237524 433304 237530 433356
rect 189902 431876 189908 431928
rect 189960 431916 189966 431928
rect 237374 431916 237380 431928
rect 189960 431888 237380 431916
rect 189960 431876 189966 431888
rect 237374 431876 237380 431888
rect 237432 431876 237438 431928
rect 198274 429156 198280 429208
rect 198332 429196 198338 429208
rect 237374 429196 237380 429208
rect 198332 429168 237380 429196
rect 198332 429156 198338 429168
rect 237374 429156 237380 429168
rect 237432 429156 237438 429208
rect 193950 427796 193956 427848
rect 194008 427836 194014 427848
rect 237374 427836 237380 427848
rect 194008 427808 237380 427836
rect 194008 427796 194014 427808
rect 237374 427796 237380 427808
rect 237432 427796 237438 427848
rect 191374 426368 191380 426420
rect 191432 426408 191438 426420
rect 237374 426408 237380 426420
rect 191432 426380 237380 426408
rect 191432 426368 191438 426380
rect 237374 426368 237380 426380
rect 237432 426368 237438 426420
rect 198366 425076 198372 425128
rect 198424 425116 198430 425128
rect 237374 425116 237380 425128
rect 198424 425088 237380 425116
rect 198424 425076 198430 425088
rect 237374 425076 237380 425088
rect 237432 425076 237438 425128
rect 191374 423648 191380 423700
rect 191432 423688 191438 423700
rect 237374 423688 237380 423700
rect 191432 423660 237380 423688
rect 191432 423648 191438 423660
rect 237374 423648 237380 423660
rect 237432 423648 237438 423700
rect 191466 422220 191472 422272
rect 191524 422260 191530 422272
rect 237374 422260 237380 422272
rect 191524 422232 237380 422260
rect 191524 422220 191530 422232
rect 237374 422220 237380 422232
rect 237432 422220 237438 422272
rect 196802 420928 196808 420980
rect 196860 420968 196866 420980
rect 237374 420968 237380 420980
rect 196860 420940 237380 420968
rect 196860 420928 196866 420940
rect 237374 420928 237380 420940
rect 237432 420928 237438 420980
rect 191466 419500 191472 419552
rect 191524 419540 191530 419552
rect 237374 419540 237380 419552
rect 191524 419512 237380 419540
rect 191524 419500 191530 419512
rect 237374 419500 237380 419512
rect 237432 419500 237438 419552
rect 501598 418140 501604 418192
rect 501656 418180 501662 418192
rect 580166 418180 580172 418192
rect 501656 418152 580172 418180
rect 501656 418140 501662 418152
rect 580166 418140 580172 418152
rect 580224 418140 580230 418192
rect 196894 415488 196900 415540
rect 196952 415528 196958 415540
rect 237466 415528 237472 415540
rect 196952 415500 237472 415528
rect 196952 415488 196958 415500
rect 237466 415488 237472 415500
rect 237524 415488 237530 415540
rect 191558 415420 191564 415472
rect 191616 415460 191622 415472
rect 237374 415460 237380 415472
rect 191616 415432 237380 415460
rect 191616 415420 191622 415432
rect 237374 415420 237380 415432
rect 237432 415420 237438 415472
rect 191282 413924 191288 413976
rect 191340 413964 191346 413976
rect 237374 413964 237380 413976
rect 191340 413936 237380 413964
rect 191340 413924 191346 413936
rect 237374 413924 237380 413936
rect 237432 413924 237438 413976
rect 196986 411272 196992 411324
rect 197044 411312 197050 411324
rect 237374 411312 237380 411324
rect 197044 411284 237380 411312
rect 197044 411272 197050 411284
rect 237374 411272 237380 411284
rect 237432 411272 237438 411324
rect 195606 407124 195612 407176
rect 195664 407164 195670 407176
rect 237374 407164 237380 407176
rect 195664 407136 237380 407164
rect 195664 407124 195670 407136
rect 237374 407124 237380 407136
rect 237432 407124 237438 407176
rect 192662 405628 192668 405680
rect 192720 405668 192726 405680
rect 237374 405668 237380 405680
rect 192720 405640 237380 405668
rect 192720 405628 192726 405640
rect 237374 405628 237380 405640
rect 237432 405628 237438 405680
rect 192846 402976 192852 403028
rect 192904 403016 192910 403028
rect 237374 403016 237380 403028
rect 192904 402988 237380 403016
rect 192904 402976 192910 402988
rect 237374 402976 237380 402988
rect 237432 402976 237438 403028
rect 188706 400120 188712 400172
rect 188764 400160 188770 400172
rect 237374 400160 237380 400172
rect 188764 400132 237380 400160
rect 188764 400120 188770 400132
rect 237374 400120 237380 400132
rect 237432 400120 237438 400172
rect 189074 398828 189080 398880
rect 189132 398868 189138 398880
rect 192662 398868 192668 398880
rect 189132 398840 192668 398868
rect 189132 398828 189138 398840
rect 192662 398828 192668 398840
rect 192720 398828 192726 398880
rect 194042 398828 194048 398880
rect 194100 398868 194106 398880
rect 237374 398868 237380 398880
rect 194100 398840 237380 398868
rect 194100 398828 194106 398840
rect 237374 398828 237380 398840
rect 237432 398828 237438 398880
rect 3326 397468 3332 397520
rect 3384 397508 3390 397520
rect 46198 397508 46204 397520
rect 3384 397480 46204 397508
rect 3384 397468 3390 397480
rect 46198 397468 46204 397480
rect 46256 397468 46262 397520
rect 189074 397468 189080 397520
rect 189132 397508 189138 397520
rect 195422 397508 195428 397520
rect 189132 397480 195428 397508
rect 189132 397468 189138 397480
rect 195422 397468 195428 397480
rect 195480 397468 195486 397520
rect 189258 396040 189264 396092
rect 189316 396080 189322 396092
rect 195514 396080 195520 396092
rect 189316 396052 195520 396080
rect 189316 396040 189322 396052
rect 195514 396040 195520 396052
rect 195572 396040 195578 396092
rect 188614 395972 188620 396024
rect 188672 396012 188678 396024
rect 237374 396012 237380 396024
rect 188672 395984 237380 396012
rect 188672 395972 188678 395984
rect 237374 395972 237380 395984
rect 237432 395972 237438 396024
rect 189074 394680 189080 394732
rect 189132 394720 189138 394732
rect 192754 394720 192760 394732
rect 189132 394692 192760 394720
rect 189132 394680 189138 394692
rect 192754 394680 192760 394692
rect 192812 394680 192818 394732
rect 194134 394680 194140 394732
rect 194192 394720 194198 394732
rect 237374 394720 237380 394732
rect 194192 394692 237380 394720
rect 194192 394680 194198 394692
rect 237374 394680 237380 394692
rect 237432 394680 237438 394732
rect 189258 393320 189264 393372
rect 189316 393360 189322 393372
rect 196710 393360 196716 393372
rect 189316 393332 196716 393360
rect 189316 393320 189322 393332
rect 196710 393320 196716 393332
rect 196768 393320 196774 393372
rect 187142 391892 187148 391944
rect 187200 391932 187206 391944
rect 237374 391932 237380 391944
rect 187200 391904 237380 391932
rect 187200 391892 187206 391904
rect 237374 391892 237380 391904
rect 237432 391892 237438 391944
rect 191282 389240 191288 389292
rect 191340 389280 191346 389292
rect 237466 389280 237472 389292
rect 191340 389252 237472 389280
rect 191340 389240 191346 389252
rect 237466 389240 237472 389252
rect 237524 389240 237530 389292
rect 189902 389172 189908 389224
rect 189960 389212 189966 389224
rect 237374 389212 237380 389224
rect 189960 389184 237380 389212
rect 189960 389172 189966 389184
rect 237374 389172 237380 389184
rect 237432 389172 237438 389224
rect 188522 387744 188528 387796
rect 188580 387784 188586 387796
rect 237374 387784 237380 387796
rect 188580 387756 237380 387784
rect 188580 387744 188586 387756
rect 237374 387744 237380 387756
rect 237432 387744 237438 387796
rect 188154 385024 188160 385076
rect 188212 385064 188218 385076
rect 237374 385064 237380 385076
rect 188212 385036 237380 385064
rect 188212 385024 188218 385036
rect 237374 385024 237380 385036
rect 237432 385024 237438 385076
rect 187050 383596 187056 383648
rect 187108 383636 187114 383648
rect 237374 383636 237380 383648
rect 187108 383608 237380 383636
rect 187108 383596 187114 383608
rect 237374 383596 237380 383608
rect 237432 383596 237438 383648
rect 186682 380876 186688 380928
rect 186740 380916 186746 380928
rect 237374 380916 237380 380928
rect 186740 380888 237380 380916
rect 186740 380876 186746 380888
rect 237374 380876 237380 380888
rect 237432 380876 237438 380928
rect 145926 379448 145932 379500
rect 145984 379488 145990 379500
rect 196802 379488 196808 379500
rect 145984 379460 196808 379488
rect 145984 379448 145990 379460
rect 196802 379448 196808 379460
rect 196860 379448 196866 379500
rect 133506 379380 133512 379432
rect 133564 379420 133570 379432
rect 194042 379420 194048 379432
rect 133564 379392 194048 379420
rect 133564 379380 133570 379392
rect 194042 379380 194048 379392
rect 194100 379380 194106 379432
rect 125962 379312 125968 379364
rect 126020 379352 126026 379364
rect 188154 379352 188160 379364
rect 126020 379324 188160 379352
rect 126020 379312 126026 379324
rect 188154 379312 188160 379324
rect 188212 379312 188218 379364
rect 128538 379244 128544 379296
rect 128596 379284 128602 379296
rect 191282 379284 191288 379296
rect 128596 379256 191288 379284
rect 128596 379244 128602 379256
rect 191282 379244 191288 379256
rect 191340 379244 191346 379296
rect 123478 379176 123484 379228
rect 123536 379216 123542 379228
rect 186682 379216 186688 379228
rect 123536 379188 186688 379216
rect 123536 379176 123542 379188
rect 186682 379176 186688 379188
rect 186740 379176 186746 379228
rect 130930 379108 130936 379160
rect 130988 379148 130994 379160
rect 194134 379148 194140 379160
rect 130988 379120 194140 379148
rect 130988 379108 130994 379120
rect 194134 379108 194140 379120
rect 194192 379108 194198 379160
rect 96430 379040 96436 379092
rect 96488 379080 96494 379092
rect 189902 379080 189908 379092
rect 96488 379052 189908 379080
rect 96488 379040 96494 379052
rect 189902 379040 189908 379052
rect 189960 379040 189966 379092
rect 102226 378972 102232 379024
rect 102284 379012 102290 379024
rect 238386 379012 238392 379024
rect 102284 378984 238392 379012
rect 102284 378972 102290 378984
rect 238386 378972 238392 378984
rect 238444 378972 238450 379024
rect 98730 378904 98736 378956
rect 98788 378944 98794 378956
rect 238570 378944 238576 378956
rect 98788 378916 238576 378944
rect 98788 378904 98794 378916
rect 238570 378904 238576 378916
rect 238628 378904 238634 378956
rect 97626 378836 97632 378888
rect 97684 378876 97690 378888
rect 238662 378876 238668 378888
rect 97684 378848 238668 378876
rect 97684 378836 97690 378848
rect 238662 378836 238668 378848
rect 238720 378836 238726 378888
rect 93946 378768 93952 378820
rect 94004 378808 94010 378820
rect 237374 378808 237380 378820
rect 94004 378780 237380 378808
rect 94004 378768 94010 378780
rect 237374 378768 237380 378780
rect 237432 378768 237438 378820
rect 148502 378700 148508 378752
rect 148560 378740 148566 378752
rect 198366 378740 198372 378752
rect 148560 378712 198372 378740
rect 148560 378700 148566 378712
rect 198366 378700 198372 378712
rect 198424 378700 198430 378752
rect 150986 378632 150992 378684
rect 151044 378672 151050 378684
rect 198274 378672 198280 378684
rect 151044 378644 198280 378672
rect 151044 378632 151050 378644
rect 198274 378632 198280 378644
rect 198332 378632 198338 378684
rect 155954 378564 155960 378616
rect 156012 378604 156018 378616
rect 198182 378604 198188 378616
rect 156012 378576 198188 378604
rect 156012 378564 156018 378576
rect 198182 378564 198188 378576
rect 198240 378564 198246 378616
rect 500310 378156 500316 378208
rect 500368 378196 500374 378208
rect 579798 378196 579804 378208
rect 500368 378168 579804 378196
rect 500368 378156 500374 378168
rect 579798 378156 579804 378168
rect 579856 378156 579862 378208
rect 47946 378088 47952 378140
rect 48004 378128 48010 378140
rect 50338 378128 50344 378140
rect 48004 378100 50344 378128
rect 48004 378088 48010 378100
rect 50338 378088 50344 378100
rect 50396 378088 50402 378140
rect 95326 378088 95332 378140
rect 95384 378128 95390 378140
rect 237466 378128 237472 378140
rect 95384 378100 237472 378128
rect 95384 378088 95390 378100
rect 237466 378088 237472 378100
rect 237524 378088 237530 378140
rect 99834 378020 99840 378072
rect 99892 378060 99898 378072
rect 238478 378060 238484 378072
rect 99892 378032 238484 378060
rect 99892 378020 99898 378032
rect 238478 378020 238484 378032
rect 238536 378020 238542 378072
rect 101306 377952 101312 378004
rect 101364 377992 101370 378004
rect 238294 377992 238300 378004
rect 101364 377964 238300 377992
rect 101364 377952 101370 377964
rect 238294 377952 238300 377964
rect 238352 377952 238358 378004
rect 103330 377884 103336 377936
rect 103388 377924 103394 377936
rect 191558 377924 191564 377936
rect 103388 377896 191564 377924
rect 103388 377884 103394 377896
rect 191558 377884 191564 377896
rect 191616 377884 191622 377936
rect 73154 377816 73160 377868
rect 73212 377856 73218 377868
rect 75178 377856 75184 377868
rect 73212 377828 75184 377856
rect 73212 377816 73218 377828
rect 75178 377816 75184 377828
rect 75236 377816 75242 377868
rect 104434 377816 104440 377868
rect 104492 377856 104498 377868
rect 191466 377856 191472 377868
rect 104492 377828 191472 377856
rect 104492 377816 104498 377828
rect 191466 377816 191472 377828
rect 191524 377816 191530 377868
rect 107562 377748 107568 377800
rect 107620 377788 107626 377800
rect 193950 377788 193956 377800
rect 107620 377760 193956 377788
rect 107620 377748 107626 377760
rect 193950 377748 193956 377760
rect 194008 377748 194014 377800
rect 105906 377680 105912 377732
rect 105964 377720 105970 377732
rect 191374 377720 191380 377732
rect 105964 377692 191380 377720
rect 105964 377680 105970 377692
rect 191374 377680 191380 377692
rect 191432 377680 191438 377732
rect 110230 377612 110236 377664
rect 110288 377652 110294 377664
rect 189810 377652 189816 377664
rect 110288 377624 189816 377652
rect 110288 377612 110294 377624
rect 189810 377612 189816 377624
rect 189868 377612 189874 377664
rect 136082 377544 136088 377596
rect 136140 377584 136146 377596
rect 192846 377584 192852 377596
rect 136140 377556 192852 377584
rect 136140 377544 136146 377556
rect 192846 377544 192852 377556
rect 192904 377544 192910 377596
rect 139026 377476 139032 377528
rect 139084 377516 139090 377528
rect 195606 377516 195612 377528
rect 139084 377488 195612 377516
rect 139084 377476 139090 377488
rect 195606 377476 195612 377488
rect 195664 377476 195670 377528
rect 120994 377408 121000 377460
rect 121052 377448 121058 377460
rect 237374 377448 237380 377460
rect 121052 377420 237380 377448
rect 121052 377408 121058 377420
rect 237374 377408 237380 377420
rect 237432 377408 237438 377460
rect 141602 377340 141608 377392
rect 141660 377380 141666 377392
rect 196986 377380 196992 377392
rect 141660 377352 196992 377380
rect 141660 377340 141666 377352
rect 196986 377340 196992 377352
rect 197044 377340 197050 377392
rect 143442 377272 143448 377324
rect 143500 377312 143506 377324
rect 196894 377312 196900 377324
rect 143500 377284 196900 377312
rect 143500 377272 143506 377284
rect 196894 377272 196900 377284
rect 196952 377272 196958 377324
rect 153378 377204 153384 377256
rect 153436 377244 153442 377256
rect 188798 377244 188804 377256
rect 153436 377216 188804 377244
rect 153436 377204 153442 377216
rect 188798 377204 188804 377216
rect 188856 377204 188862 377256
rect 78306 377000 78312 377052
rect 78364 377040 78370 377052
rect 79318 377040 79324 377052
rect 78364 377012 79324 377040
rect 78364 377000 78370 377012
rect 79318 377000 79324 377012
rect 79376 377000 79382 377052
rect 91738 377000 91744 377052
rect 91796 377040 91802 377052
rect 93118 377040 93124 377052
rect 91796 377012 93124 377040
rect 91796 377000 91802 377012
rect 93118 377000 93124 377012
rect 93176 377000 93182 377052
rect 92842 376660 92848 376712
rect 92900 376700 92906 376712
rect 237374 376700 237380 376712
rect 92900 376672 237380 376700
rect 92900 376660 92906 376672
rect 237374 376660 237380 376672
rect 237432 376660 237438 376712
rect 49326 375980 49332 376032
rect 49384 376020 49390 376032
rect 238294 376020 238300 376032
rect 49384 375992 238300 376020
rect 49384 375980 49390 375992
rect 238294 375980 238300 375992
rect 238352 375980 238358 376032
rect 118602 373940 118608 373992
rect 118660 373980 118666 373992
rect 237374 373980 237380 373992
rect 118660 373952 237380 373980
rect 118660 373940 118666 373952
rect 237374 373940 237380 373952
rect 237432 373940 237438 373992
rect 92290 372512 92296 372564
rect 92348 372552 92354 372564
rect 237374 372552 237380 372564
rect 92348 372524 237380 372552
rect 92348 372512 92354 372524
rect 237374 372512 237380 372524
rect 237432 372512 237438 372564
rect 48222 370472 48228 370524
rect 48280 370512 48286 370524
rect 148318 370512 148324 370524
rect 48280 370484 148324 370512
rect 48280 370472 48286 370484
rect 148318 370472 148324 370484
rect 148376 370472 148382 370524
rect 91002 368432 91008 368484
rect 91060 368472 91066 368484
rect 237466 368472 237472 368484
rect 91060 368444 237472 368472
rect 91060 368432 91066 368444
rect 237466 368432 237472 368444
rect 237524 368432 237530 368484
rect 117222 368364 117228 368416
rect 117280 368404 117286 368416
rect 237374 368404 237380 368416
rect 117280 368376 237380 368404
rect 117280 368364 117286 368376
rect 237374 368364 237380 368376
rect 237432 368364 237438 368416
rect 47854 367752 47860 367804
rect 47912 367792 47918 367804
rect 122098 367792 122104 367804
rect 47912 367764 122104 367792
rect 47912 367752 47918 367764
rect 122098 367752 122104 367764
rect 122156 367752 122162 367804
rect 48038 365644 48044 365696
rect 48096 365684 48102 365696
rect 50430 365684 50436 365696
rect 48096 365656 50436 365684
rect 48096 365644 48102 365656
rect 50430 365644 50436 365656
rect 50488 365644 50494 365696
rect 501690 364352 501696 364404
rect 501748 364392 501754 364404
rect 580166 364392 580172 364404
rect 501748 364364 580172 364392
rect 501748 364352 501754 364364
rect 580166 364352 580172 364364
rect 580224 364352 580230 364404
rect 89530 364284 89536 364336
rect 89588 364324 89594 364336
rect 237466 364324 237472 364336
rect 89588 364296 237472 364324
rect 89588 364284 89594 364296
rect 237466 364284 237472 364296
rect 237524 364284 237530 364336
rect 114462 364216 114468 364268
rect 114520 364256 114526 364268
rect 237374 364256 237380 364268
rect 114520 364228 237380 364256
rect 114520 364216 114526 364228
rect 237374 364216 237380 364228
rect 237432 364216 237438 364268
rect 188430 361496 188436 361548
rect 188488 361536 188494 361548
rect 237374 361536 237380 361548
rect 188488 361508 237380 361536
rect 188488 361496 188494 361508
rect 237374 361496 237380 361508
rect 237432 361496 237438 361548
rect 111702 360136 111708 360188
rect 111760 360176 111766 360188
rect 237374 360176 237380 360188
rect 111760 360148 237380 360176
rect 111760 360136 111766 360148
rect 237374 360136 237380 360148
rect 237432 360136 237438 360188
rect 48130 359456 48136 359508
rect 48188 359496 48194 359508
rect 167638 359496 167644 359508
rect 48188 359468 167644 359496
rect 48188 359456 48194 359468
rect 167638 359456 167644 359468
rect 167696 359456 167702 359508
rect 88150 358708 88156 358760
rect 88208 358748 88214 358760
rect 237374 358748 237380 358760
rect 88208 358720 237380 358748
rect 88208 358708 88214 358720
rect 237374 358708 237380 358720
rect 237432 358708 237438 358760
rect 108942 355988 108948 356040
rect 109000 356028 109006 356040
rect 237374 356028 237380 356040
rect 109000 356000 237380 356028
rect 109000 355988 109006 356000
rect 237374 355988 237380 356000
rect 237432 355988 237438 356040
rect 88242 354628 88248 354680
rect 88300 354668 88306 354680
rect 237374 354668 237380 354680
rect 88300 354640 237380 354668
rect 88300 354628 88306 354640
rect 237374 354628 237380 354640
rect 237432 354628 237438 354680
rect 106182 351840 106188 351892
rect 106240 351880 106246 351892
rect 237374 351880 237380 351892
rect 106240 351852 237380 351880
rect 106240 351840 106246 351852
rect 237374 351840 237380 351852
rect 237432 351840 237438 351892
rect 86770 350480 86776 350532
rect 86828 350520 86834 350532
rect 237374 350520 237380 350532
rect 86828 350492 237380 350520
rect 86828 350480 86834 350492
rect 237374 350480 237380 350492
rect 237432 350480 237438 350532
rect 104802 347692 104808 347744
rect 104860 347732 104866 347744
rect 237466 347732 237472 347744
rect 104860 347704 237472 347732
rect 104860 347692 104866 347704
rect 237466 347692 237472 347704
rect 237524 347692 237530 347744
rect 193858 347624 193864 347676
rect 193916 347664 193922 347676
rect 237374 347664 237380 347676
rect 193916 347636 237380 347664
rect 193916 347624 193922 347636
rect 237374 347624 237380 347636
rect 237432 347624 237438 347676
rect 49418 347012 49424 347064
rect 49476 347052 49482 347064
rect 238018 347052 238024 347064
rect 49476 347024 238024 347052
rect 49476 347012 49482 347024
rect 238018 347012 238024 347024
rect 238076 347012 238082 347064
rect 85482 346332 85488 346384
rect 85540 346372 85546 346384
rect 237374 346372 237380 346384
rect 85540 346344 237380 346372
rect 85540 346332 85546 346344
rect 237374 346332 237380 346344
rect 237432 346332 237438 346384
rect 189718 343544 189724 343596
rect 189776 343584 189782 343596
rect 237374 343584 237380 343596
rect 189776 343556 237380 343584
rect 189776 343544 189782 343556
rect 237374 343544 237380 343556
rect 237432 343544 237438 343596
rect 84010 342184 84016 342236
rect 84068 342224 84074 342236
rect 237466 342224 237472 342236
rect 84068 342196 237472 342224
rect 84068 342184 84074 342196
rect 237466 342184 237472 342196
rect 237524 342184 237530 342236
rect 102042 342116 102048 342168
rect 102100 342156 102106 342168
rect 237374 342156 237380 342168
rect 102100 342128 237380 342156
rect 102100 342116 102106 342128
rect 237374 342116 237380 342128
rect 237432 342116 237438 342168
rect 3878 340144 3884 340196
rect 3936 340184 3942 340196
rect 191190 340184 191196 340196
rect 3936 340156 191196 340184
rect 3936 340144 3942 340156
rect 191190 340144 191196 340156
rect 191248 340144 191254 340196
rect 198090 339396 198096 339448
rect 198148 339436 198154 339448
rect 237374 339436 237380 339448
rect 198148 339408 237380 339436
rect 198148 339396 198154 339408
rect 237374 339396 237380 339408
rect 237432 339396 237438 339448
rect 82722 338036 82728 338088
rect 82780 338076 82786 338088
rect 237466 338076 237472 338088
rect 82780 338048 237472 338076
rect 82780 338036 82786 338048
rect 237466 338036 237472 338048
rect 237524 338036 237530 338088
rect 99282 337968 99288 338020
rect 99340 338008 99346 338020
rect 237374 338008 237380 338020
rect 99340 337980 237380 338008
rect 99340 337968 99346 337980
rect 237374 337968 237380 337980
rect 237432 337968 237438 338020
rect 173710 336676 173716 336728
rect 173768 336716 173774 336728
rect 237374 336716 237380 336728
rect 173768 336688 237380 336716
rect 173768 336676 173774 336688
rect 237374 336676 237380 336688
rect 237432 336676 237438 336728
rect 50430 335248 50436 335300
rect 50488 335288 50494 335300
rect 237374 335288 237380 335300
rect 50488 335260 237380 335288
rect 50488 335248 50494 335260
rect 237374 335248 237380 335260
rect 237432 335248 237438 335300
rect 197998 335180 198004 335232
rect 198056 335220 198062 335232
rect 237466 335220 237472 335232
rect 198056 335192 237472 335220
rect 198056 335180 198062 335192
rect 237466 335180 237472 335192
rect 237524 335180 237530 335232
rect 96522 333888 96528 333940
rect 96580 333928 96586 333940
rect 237374 333928 237380 333940
rect 96580 333900 237380 333928
rect 96580 333888 96586 333900
rect 237374 333888 237380 333900
rect 237432 333888 237438 333940
rect 81158 332528 81164 332580
rect 81216 332568 81222 332580
rect 237374 332568 237380 332580
rect 81216 332540 237380 332568
rect 81216 332528 81222 332540
rect 237374 332528 237380 332540
rect 237432 332528 237438 332580
rect 173802 332460 173808 332512
rect 173860 332500 173866 332512
rect 237466 332500 237472 332512
rect 173860 332472 237472 332500
rect 173860 332460 173866 332472
rect 237466 332460 237472 332472
rect 237524 332460 237530 332512
rect 167638 331168 167644 331220
rect 167696 331208 167702 331220
rect 237374 331208 237380 331220
rect 167696 331180 237380 331208
rect 167696 331168 167702 331180
rect 237374 331168 237380 331180
rect 237432 331168 237438 331220
rect 93762 329740 93768 329792
rect 93820 329780 93826 329792
rect 237374 329780 237380 329792
rect 93820 329752 237380 329780
rect 93820 329740 93826 329752
rect 237374 329740 237380 329752
rect 237432 329740 237438 329792
rect 81250 328380 81256 328432
rect 81308 328420 81314 328432
rect 237374 328420 237380 328432
rect 81308 328392 237380 328420
rect 81308 328380 81314 328392
rect 237374 328380 237380 328392
rect 237432 328380 237438 328432
rect 196710 328312 196716 328364
rect 196768 328352 196774 328364
rect 237466 328352 237472 328364
rect 196768 328324 237472 328352
rect 196768 328312 196774 328324
rect 237466 328312 237472 328324
rect 237524 328312 237530 328364
rect 50338 327020 50344 327072
rect 50396 327060 50402 327072
rect 237374 327060 237380 327072
rect 50396 327032 237380 327060
rect 50396 327020 50402 327032
rect 237374 327020 237380 327032
rect 237432 327020 237438 327072
rect 93118 325592 93124 325644
rect 93176 325632 93182 325644
rect 237374 325632 237380 325644
rect 93176 325604 237380 325632
rect 93176 325592 93182 325604
rect 237374 325592 237380 325604
rect 237432 325592 237438 325644
rect 235350 325524 235356 325576
rect 235408 325564 235414 325576
rect 237466 325564 237472 325576
rect 235408 325536 237472 325564
rect 235408 325524 235414 325536
rect 237466 325524 237472 325536
rect 237524 325524 237530 325576
rect 499022 324300 499028 324352
rect 499080 324340 499086 324352
rect 579982 324340 579988 324352
rect 499080 324312 579988 324340
rect 499080 324300 499086 324312
rect 579982 324300 579988 324312
rect 580040 324300 580046 324352
rect 79962 324232 79968 324284
rect 80020 324272 80026 324284
rect 237374 324272 237380 324284
rect 80020 324244 237380 324272
rect 80020 324232 80026 324244
rect 237374 324232 237380 324244
rect 237432 324232 237438 324284
rect 192754 322872 192760 322924
rect 192812 322912 192818 322924
rect 237374 322912 237380 322924
rect 192812 322884 237380 322912
rect 192812 322872 192818 322884
rect 237374 322872 237380 322884
rect 237432 322872 237438 322924
rect 235258 321512 235264 321564
rect 235316 321552 235322 321564
rect 237374 321552 237380 321564
rect 235316 321524 237380 321552
rect 235316 321512 235322 321524
rect 237374 321512 237380 321524
rect 237432 321512 237438 321564
rect 78490 320084 78496 320136
rect 78548 320124 78554 320136
rect 237466 320124 237472 320136
rect 78548 320096 237472 320124
rect 78548 320084 78554 320096
rect 237466 320084 237472 320096
rect 237524 320084 237530 320136
rect 89622 320016 89628 320068
rect 89680 320056 89686 320068
rect 237374 320056 237380 320068
rect 89680 320028 237380 320056
rect 89680 320016 89686 320028
rect 237374 320016 237380 320028
rect 237432 320016 237438 320068
rect 195514 318724 195520 318776
rect 195572 318764 195578 318776
rect 237374 318764 237380 318776
rect 195572 318736 237380 318764
rect 195572 318724 195578 318736
rect 237374 318724 237380 318736
rect 237432 318724 237438 318776
rect 73062 317364 73068 317416
rect 73120 317404 73126 317416
rect 237374 317404 237380 317416
rect 73120 317376 237380 317404
rect 73120 317364 73126 317376
rect 237374 317364 237380 317376
rect 237432 317364 237438 317416
rect 86862 315936 86868 315988
rect 86920 315976 86926 315988
rect 237374 315976 237380 315988
rect 86920 315948 237380 315976
rect 86920 315936 86926 315948
rect 237374 315936 237380 315948
rect 237432 315936 237438 315988
rect 77202 314576 77208 314628
rect 77260 314616 77266 314628
rect 237374 314616 237380 314628
rect 77260 314588 237380 314616
rect 77260 314576 77266 314588
rect 237374 314576 237380 314588
rect 237432 314576 237438 314628
rect 49234 313216 49240 313268
rect 49292 313256 49298 313268
rect 237466 313256 237472 313268
rect 49292 313228 237472 313256
rect 49292 313216 49298 313228
rect 237466 313216 237472 313228
rect 237524 313216 237530 313268
rect 195422 313148 195428 313200
rect 195480 313188 195486 313200
rect 237374 313188 237380 313200
rect 195480 313160 237380 313188
rect 195480 313148 195486 313160
rect 237374 313148 237380 313160
rect 237432 313148 237438 313200
rect 71682 311788 71688 311840
rect 71740 311828 71746 311840
rect 237374 311828 237380 311840
rect 71740 311800 237380 311828
rect 71740 311788 71746 311800
rect 237374 311788 237380 311800
rect 237432 311788 237438 311840
rect 84102 310428 84108 310480
rect 84160 310468 84166 310480
rect 237466 310468 237472 310480
rect 84160 310440 237472 310468
rect 84160 310428 84166 310440
rect 237466 310428 237472 310440
rect 237524 310428 237530 310480
rect 196618 310360 196624 310412
rect 196676 310400 196682 310412
rect 237374 310400 237380 310412
rect 196676 310372 237380 310400
rect 196676 310360 196682 310372
rect 237374 310360 237380 310372
rect 237432 310360 237438 310412
rect 75822 309068 75828 309120
rect 75880 309108 75886 309120
rect 237374 309108 237380 309120
rect 75880 309080 237380 309108
rect 75880 309068 75886 309080
rect 237374 309068 237380 309080
rect 237432 309068 237438 309120
rect 192662 309000 192668 309052
rect 192720 309040 192726 309052
rect 237466 309040 237472 309052
rect 192720 309012 237472 309040
rect 192720 309000 192726 309012
rect 237466 309000 237472 309012
rect 237524 309000 237530 309052
rect 49602 307708 49608 307760
rect 49660 307748 49666 307760
rect 237374 307748 237380 307760
rect 49660 307720 237380 307748
rect 49660 307708 49666 307720
rect 237374 307708 237380 307720
rect 237432 307708 237438 307760
rect 70302 306280 70308 306332
rect 70360 306320 70366 306332
rect 237374 306320 237380 306332
rect 70360 306292 237380 306320
rect 70360 306280 70366 306292
rect 237374 306280 237380 306292
rect 237432 306280 237438 306332
rect 188338 306212 188344 306264
rect 188396 306252 188402 306264
rect 237466 306252 237472 306264
rect 188396 306224 237472 306252
rect 188396 306212 188402 306224
rect 237466 306212 237472 306224
rect 237524 306212 237530 306264
rect 3142 304988 3148 305040
rect 3200 305028 3206 305040
rect 228358 305028 228364 305040
rect 3200 305000 228364 305028
rect 3200 304988 3206 305000
rect 228358 304988 228364 305000
rect 228416 304988 228422 305040
rect 81342 304920 81348 304972
rect 81400 304960 81406 304972
rect 237374 304960 237380 304972
rect 81400 304932 237380 304960
rect 81400 304920 81406 304932
rect 237374 304920 237380 304932
rect 237432 304920 237438 304972
rect 74350 303560 74356 303612
rect 74408 303600 74414 303612
rect 237374 303600 237380 303612
rect 74408 303572 237380 303600
rect 74408 303560 74414 303572
rect 237374 303560 237380 303572
rect 237432 303560 237438 303612
rect 192570 303492 192576 303544
rect 192628 303532 192634 303544
rect 237466 303532 237472 303544
rect 192628 303504 237472 303532
rect 192628 303492 192634 303504
rect 237466 303492 237472 303504
rect 237524 303492 237530 303544
rect 67542 302132 67548 302184
rect 67600 302172 67606 302184
rect 237374 302172 237380 302184
rect 67600 302144 237380 302172
rect 67600 302132 67606 302144
rect 237374 302132 237380 302144
rect 237432 302132 237438 302184
rect 68922 300772 68928 300824
rect 68980 300812 68986 300824
rect 237374 300812 237380 300824
rect 68980 300784 237380 300812
rect 68980 300772 68986 300784
rect 237374 300772 237380 300784
rect 237432 300772 237438 300824
rect 195238 300704 195244 300756
rect 195296 300744 195302 300756
rect 237466 300744 237472 300756
rect 195296 300716 237472 300744
rect 195296 300704 195302 300716
rect 237466 300704 237472 300716
rect 237524 300704 237530 300756
rect 75178 299412 75184 299464
rect 75236 299452 75242 299464
rect 237466 299452 237472 299464
rect 75236 299424 237472 299452
rect 75236 299412 75242 299424
rect 237466 299412 237472 299424
rect 237524 299412 237530 299464
rect 79318 299344 79324 299396
rect 79376 299384 79382 299396
rect 237374 299384 237380 299396
rect 79376 299356 237380 299384
rect 79376 299344 79382 299356
rect 237374 299344 237380 299356
rect 237432 299344 237438 299396
rect 192478 298052 192484 298104
rect 192536 298092 192542 298104
rect 237374 298092 237380 298104
rect 192536 298064 237380 298092
rect 192536 298052 192542 298064
rect 237374 298052 237380 298064
rect 237432 298052 237438 298104
rect 66162 296624 66168 296676
rect 66220 296664 66226 296676
rect 237374 296664 237380 296676
rect 66220 296636 237380 296664
rect 66220 296624 66226 296636
rect 237374 296624 237380 296636
rect 237432 296624 237438 296676
rect 148318 296556 148324 296608
rect 148376 296596 148382 296608
rect 237466 296596 237472 296608
rect 148376 296568 237472 296596
rect 148376 296556 148382 296568
rect 237466 296556 237472 296568
rect 237524 296556 237530 296608
rect 195330 295264 195336 295316
rect 195388 295304 195394 295316
rect 237374 295304 237380 295316
rect 195388 295276 237380 295304
rect 195388 295264 195394 295276
rect 237374 295264 237380 295276
rect 237432 295264 237438 295316
rect 122098 293904 122104 293956
rect 122156 293944 122162 293956
rect 237374 293944 237380 293956
rect 122156 293916 237380 293944
rect 122156 293904 122162 293916
rect 237374 293904 237380 293916
rect 237432 293904 237438 293956
rect 157242 292612 157248 292664
rect 157300 292652 157306 292664
rect 237374 292652 237380 292664
rect 157300 292624 237380 292652
rect 157300 292612 157306 292624
rect 237374 292612 237380 292624
rect 237432 292612 237438 292664
rect 3326 292544 3332 292596
rect 3384 292584 3390 292596
rect 236638 292584 236644 292596
rect 3384 292556 236644 292584
rect 3384 292544 3390 292556
rect 236638 292544 236644 292556
rect 236696 292544 236702 292596
rect 235258 291184 235264 291236
rect 235316 291224 235322 291236
rect 237374 291224 237380 291236
rect 235316 291196 237380 291224
rect 235316 291184 235322 291196
rect 237374 291184 237380 291196
rect 237432 291184 237438 291236
rect 154482 289824 154488 289876
rect 154540 289864 154546 289876
rect 237374 289864 237380 289876
rect 154540 289836 237380 289864
rect 154540 289824 154546 289836
rect 237374 289824 237380 289836
rect 237432 289824 237438 289876
rect 235350 288464 235356 288516
rect 235408 288504 235414 288516
rect 237466 288504 237472 288516
rect 235408 288476 237472 288504
rect 235408 288464 235414 288476
rect 237466 288464 237472 288476
rect 237524 288464 237530 288516
rect 235442 288396 235448 288448
rect 235500 288436 235506 288448
rect 237374 288436 237380 288448
rect 235500 288408 237380 288436
rect 235500 288396 235506 288408
rect 237374 288396 237380 288408
rect 237432 288396 237438 288448
rect 151722 287036 151728 287088
rect 151780 287076 151786 287088
rect 237374 287076 237380 287088
rect 151780 287048 237380 287076
rect 151780 287036 151786 287048
rect 237374 287036 237380 287048
rect 237432 287036 237438 287088
rect 170674 286560 170680 286612
rect 170732 286600 170738 286612
rect 192478 286600 192484 286612
rect 170732 286572 192484 286600
rect 170732 286560 170738 286572
rect 192478 286560 192484 286572
rect 192536 286560 192542 286612
rect 169662 286492 169668 286544
rect 169720 286532 169726 286544
rect 192570 286532 192576 286544
rect 169720 286504 192576 286532
rect 169720 286492 169726 286504
rect 192570 286492 192576 286504
rect 192628 286492 192634 286544
rect 144822 286424 144828 286476
rect 144880 286464 144886 286476
rect 186774 286464 186780 286476
rect 144880 286436 186780 286464
rect 144880 286424 144886 286436
rect 186774 286424 186780 286436
rect 186832 286424 186838 286476
rect 141878 286356 141884 286408
rect 141936 286396 141942 286408
rect 187326 286396 187332 286408
rect 141936 286368 187332 286396
rect 141936 286356 141942 286368
rect 187326 286356 187332 286368
rect 187384 286356 187390 286408
rect 139302 286288 139308 286340
rect 139360 286328 139366 286340
rect 187234 286328 187240 286340
rect 139360 286300 187240 286328
rect 139360 286288 139366 286300
rect 187234 286288 187240 286300
rect 187292 286288 187298 286340
rect 136542 286220 136548 286272
rect 136600 286260 136606 286272
rect 187142 286260 187148 286272
rect 136600 286232 187148 286260
rect 136600 286220 136606 286232
rect 187142 286220 187148 286232
rect 187200 286220 187206 286272
rect 126882 286152 126888 286204
rect 126940 286192 126946 286204
rect 187050 286192 187056 286204
rect 126940 286164 187056 286192
rect 126940 286152 126946 286164
rect 187050 286152 187056 286164
rect 187108 286152 187114 286204
rect 124122 286084 124128 286136
rect 124180 286124 124186 286136
rect 186958 286124 186964 286136
rect 124180 286096 186964 286124
rect 124180 286084 124186 286096
rect 186958 286084 186964 286096
rect 187016 286084 187022 286136
rect 108942 286016 108948 286068
rect 109000 286056 109006 286068
rect 194042 286056 194048 286068
rect 109000 286028 194048 286056
rect 109000 286016 109006 286028
rect 194042 286016 194048 286028
rect 194100 286016 194106 286068
rect 106182 285948 106188 286000
rect 106240 285988 106246 286000
rect 191466 285988 191472 286000
rect 106240 285960 191472 285988
rect 106240 285948 106246 285960
rect 191466 285948 191472 285960
rect 191524 285948 191530 286000
rect 104802 285880 104808 285932
rect 104860 285920 104866 285932
rect 192754 285920 192760 285932
rect 104860 285892 192760 285920
rect 104860 285880 104866 285892
rect 192754 285880 192760 285892
rect 192812 285880 192818 285932
rect 238110 285920 238116 285932
rect 219406 285892 238116 285920
rect 118602 285812 118608 285864
rect 118660 285852 118666 285864
rect 219406 285852 219434 285892
rect 238110 285880 238116 285892
rect 238168 285880 238174 285932
rect 238202 285852 238208 285864
rect 118660 285824 219434 285852
rect 233620 285824 238208 285852
rect 118660 285812 118666 285824
rect 114462 285744 114468 285796
rect 114520 285784 114526 285796
rect 233620 285784 233648 285824
rect 238202 285812 238208 285824
rect 238260 285812 238266 285864
rect 114520 285756 233648 285784
rect 114520 285744 114526 285756
rect 235534 285744 235540 285796
rect 235592 285784 235598 285796
rect 237466 285784 237472 285796
rect 235592 285756 237472 285784
rect 235592 285744 235598 285756
rect 237466 285744 237472 285756
rect 237524 285744 237530 285796
rect 83734 285676 83740 285728
rect 83792 285716 83798 285728
rect 232590 285716 232596 285728
rect 83792 285688 232596 285716
rect 83792 285676 83798 285688
rect 232590 285676 232596 285688
rect 232648 285676 232654 285728
rect 235626 285676 235632 285728
rect 235684 285716 235690 285728
rect 237374 285716 237380 285728
rect 235684 285688 237380 285716
rect 235684 285676 235690 285688
rect 237374 285676 237380 285688
rect 237432 285676 237438 285728
rect 92382 285608 92388 285660
rect 92440 285648 92446 285660
rect 191282 285648 191288 285660
rect 92440 285620 191288 285648
rect 92440 285608 92446 285620
rect 191282 285608 191288 285620
rect 191340 285608 191346 285660
rect 93670 285540 93676 285592
rect 93728 285580 93734 285592
rect 195238 285580 195244 285592
rect 93728 285552 195244 285580
rect 93728 285540 93734 285552
rect 195238 285540 195244 285552
rect 195296 285540 195302 285592
rect 96522 285472 96528 285524
rect 96580 285512 96586 285524
rect 198090 285512 198096 285524
rect 96580 285484 198096 285512
rect 96580 285472 96586 285484
rect 198090 285472 198096 285484
rect 198148 285472 198154 285524
rect 86862 285404 86868 285456
rect 86920 285444 86926 285456
rect 189718 285444 189724 285456
rect 86920 285416 189724 285444
rect 86920 285404 86926 285416
rect 189718 285404 189724 285416
rect 189776 285404 189782 285456
rect 133782 285336 133788 285388
rect 133840 285376 133846 285388
rect 237834 285376 237840 285388
rect 133840 285348 237840 285376
rect 133840 285336 133846 285348
rect 237834 285336 237840 285348
rect 237892 285336 237898 285388
rect 89622 285268 89628 285320
rect 89680 285308 89686 285320
rect 193858 285308 193864 285320
rect 89680 285280 193864 285308
rect 89680 285268 89686 285280
rect 193858 285268 193864 285280
rect 193916 285268 193922 285320
rect 131114 285200 131120 285252
rect 131172 285240 131178 285252
rect 238478 285240 238484 285252
rect 131172 285212 238484 285240
rect 131172 285200 131178 285212
rect 238478 285200 238484 285212
rect 238536 285200 238542 285252
rect 128722 285132 128728 285184
rect 128780 285172 128786 285184
rect 238662 285172 238668 285184
rect 128780 285144 238668 285172
rect 128780 285132 128786 285144
rect 238662 285132 238668 285144
rect 238720 285132 238726 285184
rect 116210 285064 116216 285116
rect 116268 285104 116274 285116
rect 238570 285104 238576 285116
rect 116268 285076 238576 285104
rect 116268 285064 116274 285076
rect 238570 285064 238576 285076
rect 238628 285064 238634 285116
rect 111058 284996 111064 285048
rect 111116 285036 111122 285048
rect 238386 285036 238392 285048
rect 111116 285008 238392 285036
rect 111116 284996 111122 285008
rect 238386 284996 238392 285008
rect 238444 284996 238450 285048
rect 98546 284928 98552 284980
rect 98604 284968 98610 284980
rect 238018 284968 238024 284980
rect 98604 284940 238024 284968
rect 98604 284928 98610 284940
rect 238018 284928 238024 284940
rect 238076 284928 238082 284980
rect 148594 284860 148600 284912
rect 148652 284900 148658 284912
rect 237374 284900 237380 284912
rect 148652 284872 237380 284900
rect 148652 284860 148658 284872
rect 237374 284860 237380 284872
rect 237432 284860 237438 284912
rect 101306 284792 101312 284844
rect 101364 284832 101370 284844
rect 189902 284832 189908 284844
rect 101364 284804 189908 284832
rect 101364 284792 101370 284804
rect 189902 284792 189908 284804
rect 189960 284792 189966 284844
rect 146018 284724 146024 284776
rect 146076 284764 146082 284776
rect 186682 284764 186688 284776
rect 146076 284736 186688 284764
rect 146076 284724 146082 284736
rect 186682 284724 186688 284736
rect 186740 284724 186746 284776
rect 235810 282956 235816 283008
rect 235868 282996 235874 283008
rect 237374 282996 237380 283008
rect 235868 282968 237380 282996
rect 235868 282956 235874 282968
rect 237374 282956 237380 282968
rect 237432 282956 237438 283008
rect 235718 282888 235724 282940
rect 235776 282928 235782 282940
rect 237466 282928 237472 282940
rect 235776 282900 237472 282928
rect 235776 282888 235782 282900
rect 237466 282888 237472 282900
rect 237524 282888 237530 282940
rect 186682 282820 186688 282872
rect 186740 282860 186746 282872
rect 237374 282860 237380 282872
rect 186740 282832 237380 282860
rect 186740 282820 186746 282832
rect 237374 282820 237380 282832
rect 237432 282820 237438 282872
rect 192662 280236 192668 280288
rect 192720 280276 192726 280288
rect 237374 280276 237380 280288
rect 192720 280248 237380 280276
rect 192720 280236 192726 280248
rect 237374 280236 237380 280248
rect 237432 280236 237438 280288
rect 187602 280168 187608 280220
rect 187660 280208 187666 280220
rect 237466 280208 237472 280220
rect 187660 280180 237472 280208
rect 187660 280168 187666 280180
rect 237466 280168 237472 280180
rect 237524 280168 237530 280220
rect 186774 280100 186780 280152
rect 186832 280140 186838 280152
rect 237374 280140 237380 280152
rect 186832 280112 237380 280140
rect 186832 280100 186838 280112
rect 237374 280100 237380 280112
rect 237432 280100 237438 280152
rect 189994 278740 190000 278792
rect 190052 278780 190058 278792
rect 215938 278780 215944 278792
rect 190052 278752 215944 278780
rect 190052 278740 190058 278752
rect 215938 278740 215944 278752
rect 215996 278740 216002 278792
rect 187326 277312 187332 277364
rect 187384 277352 187390 277364
rect 237374 277352 237380 277364
rect 187384 277324 237380 277352
rect 187384 277312 187390 277324
rect 237374 277312 237380 277324
rect 237432 277312 237438 277364
rect 189810 274660 189816 274712
rect 189868 274700 189874 274712
rect 237466 274700 237472 274712
rect 189868 274672 237472 274700
rect 189868 274660 189874 274672
rect 237466 274660 237472 274672
rect 237524 274660 237530 274712
rect 187234 274592 187240 274644
rect 187292 274632 187298 274644
rect 237374 274632 237380 274644
rect 187292 274604 237380 274632
rect 187292 274592 187298 274604
rect 237374 274592 237380 274604
rect 237432 274592 237438 274644
rect 499022 271872 499028 271924
rect 499080 271912 499086 271924
rect 579798 271912 579804 271924
rect 499080 271884 579804 271912
rect 499080 271872 499086 271884
rect 579798 271872 579804 271884
rect 579856 271872 579862 271924
rect 187142 271804 187148 271856
rect 187200 271844 187206 271856
rect 237374 271844 237380 271856
rect 187200 271816 237380 271844
rect 187200 271804 187206 271816
rect 237374 271804 237380 271816
rect 237432 271804 237438 271856
rect 197998 267724 198004 267776
rect 198056 267764 198062 267776
rect 237374 267764 237380 267776
rect 198056 267736 237380 267764
rect 198056 267724 198062 267736
rect 237374 267724 237380 267736
rect 237432 267724 237438 267776
rect 188338 262216 188344 262268
rect 188396 262256 188402 262268
rect 237374 262256 237380 262268
rect 188396 262228 237380 262256
rect 188396 262216 188402 262228
rect 237374 262216 237380 262228
rect 237432 262216 237438 262268
rect 187050 262148 187056 262200
rect 187108 262188 187114 262200
rect 237466 262188 237472 262200
rect 187108 262160 237472 262188
rect 187108 262148 187114 262160
rect 237466 262148 237472 262160
rect 237524 262148 237530 262200
rect 187142 260856 187148 260908
rect 187200 260896 187206 260908
rect 237374 260896 237380 260908
rect 187200 260868 237380 260896
rect 187200 260856 187206 260868
rect 237374 260856 237380 260868
rect 237432 260856 237438 260908
rect 196618 259496 196624 259548
rect 196676 259536 196682 259548
rect 237374 259536 237380 259548
rect 196676 259508 237380 259536
rect 196676 259496 196682 259508
rect 237374 259496 237380 259508
rect 237432 259496 237438 259548
rect 187326 259428 187332 259480
rect 187384 259468 187390 259480
rect 237466 259468 237472 259480
rect 187384 259440 237472 259468
rect 187384 259428 187390 259440
rect 237466 259428 237472 259440
rect 237524 259428 237530 259480
rect 186958 259360 186964 259412
rect 187016 259400 187022 259412
rect 237374 259400 237380 259412
rect 187016 259372 237380 259400
rect 187016 259360 187022 259372
rect 237374 259360 237380 259372
rect 237432 259360 237438 259412
rect 500402 258068 500408 258120
rect 500460 258108 500466 258120
rect 579982 258108 579988 258120
rect 500460 258080 579988 258108
rect 500460 258068 500466 258080
rect 579982 258068 579988 258080
rect 580040 258068 580046 258120
rect 235902 256776 235908 256828
rect 235960 256816 235966 256828
rect 237466 256816 237472 256828
rect 235960 256788 237472 256816
rect 235960 256776 235966 256788
rect 237466 256776 237472 256788
rect 237524 256776 237530 256828
rect 188430 256708 188436 256760
rect 188488 256748 188494 256760
rect 237374 256748 237380 256760
rect 188488 256720 237380 256748
rect 188488 256708 188494 256720
rect 237374 256708 237380 256720
rect 237432 256708 237438 256760
rect 2774 254056 2780 254108
rect 2832 254096 2838 254108
rect 4798 254096 4804 254108
rect 2832 254068 4804 254096
rect 2832 254056 2838 254068
rect 4798 254056 4804 254068
rect 4856 254056 4862 254108
rect 196710 253988 196716 254040
rect 196768 254028 196774 254040
rect 237466 254028 237472 254040
rect 196768 254000 237472 254028
rect 196768 253988 196774 254000
rect 237466 253988 237472 254000
rect 237524 253988 237530 254040
rect 191374 253920 191380 253972
rect 191432 253960 191438 253972
rect 237374 253960 237380 253972
rect 191432 253932 237380 253960
rect 191432 253920 191438 253932
rect 237374 253920 237380 253932
rect 237432 253920 237438 253972
rect 195330 251200 195336 251252
rect 195388 251240 195394 251252
rect 237374 251240 237380 251252
rect 195388 251212 237380 251240
rect 195388 251200 195394 251212
rect 237374 251200 237380 251212
rect 237432 251200 237438 251252
rect 195422 249772 195428 249824
rect 195480 249812 195486 249824
rect 237374 249812 237380 249824
rect 195480 249784 237380 249812
rect 195480 249772 195486 249784
rect 237374 249772 237380 249784
rect 237432 249772 237438 249824
rect 189994 248412 190000 248464
rect 190052 248452 190058 248464
rect 237374 248452 237380 248464
rect 190052 248424 237380 248452
rect 190052 248412 190058 248424
rect 237374 248412 237380 248424
rect 237432 248412 237438 248464
rect 195514 247052 195520 247104
rect 195572 247092 195578 247104
rect 237374 247092 237380 247104
rect 195572 247064 237380 247092
rect 195572 247052 195578 247064
rect 237374 247052 237380 247064
rect 237432 247052 237438 247104
rect 193950 244264 193956 244316
rect 194008 244304 194014 244316
rect 237374 244304 237380 244316
rect 194008 244276 237380 244304
rect 194008 244264 194014 244276
rect 237374 244264 237380 244276
rect 237432 244264 237438 244316
rect 194042 242836 194048 242888
rect 194100 242876 194106 242888
rect 237374 242876 237380 242888
rect 194100 242848 237380 242876
rect 194100 242836 194106 242848
rect 237374 242836 237380 242848
rect 237432 242836 237438 242888
rect 186958 241476 186964 241528
rect 187016 241516 187022 241528
rect 237374 241516 237380 241528
rect 187016 241488 237380 241516
rect 187016 241476 187022 241488
rect 237374 241476 237380 241488
rect 237432 241476 237438 241528
rect 3142 240320 3148 240372
rect 3200 240360 3206 240372
rect 6178 240360 6184 240372
rect 3200 240332 6184 240360
rect 3200 240320 3206 240332
rect 6178 240320 6184 240332
rect 6236 240320 6242 240372
rect 191558 240116 191564 240168
rect 191616 240156 191622 240168
rect 237374 240156 237380 240168
rect 191616 240128 237380 240156
rect 191616 240116 191622 240128
rect 237374 240116 237380 240128
rect 237432 240116 237438 240168
rect 191466 238688 191472 238740
rect 191524 238728 191530 238740
rect 237374 238728 237380 238740
rect 191524 238700 237380 238728
rect 191524 238688 191530 238700
rect 237374 238688 237380 238700
rect 237432 238688 237438 238740
rect 195606 235968 195612 236020
rect 195664 236008 195670 236020
rect 237374 236008 237380 236020
rect 195664 235980 237380 236008
rect 195664 235968 195670 235980
rect 237374 235968 237380 235980
rect 237432 235968 237438 236020
rect 192754 234540 192760 234592
rect 192812 234580 192818 234592
rect 237374 234580 237380 234592
rect 192812 234552 237380 234580
rect 192812 234540 192818 234552
rect 237374 234540 237380 234552
rect 237432 234540 237438 234592
rect 188522 231820 188528 231872
rect 188580 231860 188586 231872
rect 237374 231860 237380 231872
rect 188580 231832 237380 231860
rect 188580 231820 188586 231832
rect 237374 231820 237380 231832
rect 237432 231820 237438 231872
rect 189902 230392 189908 230444
rect 189960 230432 189966 230444
rect 237374 230432 237380 230444
rect 189960 230404 237380 230432
rect 189960 230392 189966 230404
rect 237374 230392 237380 230404
rect 237432 230392 237438 230444
rect 188614 227808 188620 227860
rect 188672 227848 188678 227860
rect 237466 227848 237472 227860
rect 188672 227820 237472 227848
rect 188672 227808 188678 227820
rect 237466 227808 237472 227820
rect 237524 227808 237530 227860
rect 187050 227740 187056 227792
rect 187108 227780 187114 227792
rect 237374 227780 237380 227792
rect 187108 227752 237380 227780
rect 187108 227740 187114 227752
rect 237374 227740 237380 227752
rect 237432 227740 237438 227792
rect 188706 223592 188712 223644
rect 188764 223632 188770 223644
rect 237374 223632 237380 223644
rect 188764 223604 237380 223632
rect 188764 223592 188770 223604
rect 237374 223592 237380 223604
rect 237432 223592 237438 223644
rect 194042 222232 194048 222284
rect 194100 222272 194106 222284
rect 237374 222272 237380 222284
rect 194100 222244 237380 222272
rect 194100 222232 194106 222244
rect 237374 222232 237380 222244
rect 237432 222232 237438 222284
rect 187234 222164 187240 222216
rect 187292 222204 187298 222216
rect 237466 222204 237472 222216
rect 187292 222176 237472 222204
rect 187292 222164 187298 222176
rect 237466 222164 237472 222176
rect 237524 222164 237530 222216
rect 198090 222096 198096 222148
rect 198148 222136 198154 222148
rect 237374 222136 237380 222148
rect 198148 222108 237380 222136
rect 198148 222096 198154 222108
rect 237374 222096 237380 222108
rect 237432 222096 237438 222148
rect 188890 221484 188896 221536
rect 188948 221524 188954 221536
rect 238294 221524 238300 221536
rect 188948 221496 238300 221524
rect 188948 221484 188954 221496
rect 238294 221484 238300 221496
rect 238352 221484 238358 221536
rect 188798 221416 188804 221468
rect 188856 221456 188862 221468
rect 238478 221456 238484 221468
rect 188856 221428 238484 221456
rect 188856 221416 188862 221428
rect 238478 221416 238484 221428
rect 238536 221416 238542 221468
rect 235166 220804 235172 220856
rect 235224 220844 235230 220856
rect 237466 220844 237472 220856
rect 235224 220816 237472 220844
rect 235224 220804 235230 220816
rect 237466 220804 237472 220816
rect 237524 220804 237530 220856
rect 188982 219444 188988 219496
rect 189040 219484 189046 219496
rect 237374 219484 237380 219496
rect 189040 219456 237380 219484
rect 189040 219444 189046 219456
rect 237374 219444 237380 219456
rect 237432 219444 237438 219496
rect 189074 218152 189080 218204
rect 189132 218192 189138 218204
rect 198090 218192 198096 218204
rect 189132 218164 198096 218192
rect 189132 218152 189138 218164
rect 198090 218152 198096 218164
rect 198148 218152 198154 218204
rect 192754 218084 192760 218136
rect 192812 218124 192818 218136
rect 237374 218124 237380 218136
rect 192812 218096 237380 218124
rect 192812 218084 192818 218096
rect 237374 218084 237380 218096
rect 237432 218084 237438 218136
rect 187418 218016 187424 218068
rect 187476 218056 187482 218068
rect 237466 218056 237472 218068
rect 187476 218028 237472 218056
rect 187476 218016 187482 218028
rect 237466 218016 237472 218028
rect 237524 218016 237530 218068
rect 500494 218016 500500 218068
rect 500552 218056 500558 218068
rect 579798 218056 579804 218068
rect 500552 218028 579804 218056
rect 500552 218016 500558 218028
rect 579798 218016 579804 218028
rect 579856 218016 579862 218068
rect 195238 216588 195244 216640
rect 195296 216628 195302 216640
rect 237374 216628 237380 216640
rect 195296 216600 237380 216628
rect 195296 216588 195302 216600
rect 237374 216588 237380 216600
rect 237432 216588 237438 216640
rect 189074 215296 189080 215348
rect 189132 215336 189138 215348
rect 191466 215336 191472 215348
rect 189132 215308 191472 215336
rect 189132 215296 189138 215308
rect 191466 215296 191472 215308
rect 191524 215296 191530 215348
rect 190086 213936 190092 213988
rect 190144 213976 190150 213988
rect 191650 213976 191656 213988
rect 190144 213948 191656 213976
rect 190144 213936 190150 213948
rect 191650 213936 191656 213948
rect 191708 213936 191714 213988
rect 190270 213188 190276 213240
rect 190328 213228 190334 213240
rect 237374 213228 237380 213240
rect 190328 213200 237380 213228
rect 190328 213188 190334 213200
rect 237374 213188 237380 213200
rect 237432 213188 237438 213240
rect 234982 212508 234988 212560
rect 235040 212548 235046 212560
rect 237466 212548 237472 212560
rect 235040 212520 237472 212548
rect 235040 212508 235046 212520
rect 237466 212508 237472 212520
rect 237524 212508 237530 212560
rect 191282 212440 191288 212492
rect 191340 212480 191346 212492
rect 237374 212480 237380 212492
rect 191340 212452 237380 212480
rect 191340 212440 191346 212452
rect 237374 212440 237380 212452
rect 237432 212440 237438 212492
rect 228450 209788 228456 209840
rect 228508 209828 228514 209840
rect 237466 209828 237472 209840
rect 228508 209800 237472 209828
rect 228508 209788 228514 209800
rect 237466 209788 237472 209800
rect 237524 209788 237530 209840
rect 191650 209720 191656 209772
rect 191708 209760 191714 209772
rect 237374 209760 237380 209772
rect 191708 209732 237380 209760
rect 191708 209720 191714 209732
rect 237374 209720 237380 209732
rect 237432 209720 237438 209772
rect 191282 208360 191288 208412
rect 191340 208400 191346 208412
rect 237374 208400 237380 208412
rect 191340 208372 237380 208400
rect 191340 208360 191346 208372
rect 237374 208360 237380 208372
rect 237432 208360 237438 208412
rect 193858 208292 193864 208344
rect 193916 208332 193922 208344
rect 237466 208332 237472 208344
rect 193916 208304 237472 208332
rect 193916 208292 193922 208304
rect 237466 208292 237472 208304
rect 237524 208292 237530 208344
rect 47578 207680 47584 207732
rect 47636 207720 47642 207732
rect 48222 207720 48228 207732
rect 47636 207692 48228 207720
rect 47636 207680 47642 207692
rect 48222 207680 48228 207692
rect 48280 207720 48286 207732
rect 49602 207720 49608 207732
rect 48280 207692 49608 207720
rect 48280 207680 48286 207692
rect 49602 207680 49608 207692
rect 49660 207680 49666 207732
rect 187510 205640 187516 205692
rect 187568 205680 187574 205692
rect 237466 205680 237472 205692
rect 187568 205652 237472 205680
rect 187568 205640 187574 205652
rect 237466 205640 237472 205652
rect 237524 205640 237530 205692
rect 191466 205572 191472 205624
rect 191524 205612 191530 205624
rect 237374 205612 237380 205624
rect 191524 205584 237380 205612
rect 191524 205572 191530 205584
rect 237374 205572 237380 205584
rect 237432 205572 237438 205624
rect 191466 202920 191472 202972
rect 191524 202960 191530 202972
rect 237374 202960 237380 202972
rect 191524 202932 237380 202960
rect 191524 202920 191530 202932
rect 237374 202920 237380 202932
rect 237432 202920 237438 202972
rect 188246 202852 188252 202904
rect 188304 202892 188310 202904
rect 237466 202892 237472 202904
rect 188304 202864 237472 202892
rect 188304 202852 188310 202864
rect 237466 202852 237472 202864
rect 237524 202852 237530 202904
rect 189718 202784 189724 202836
rect 189776 202824 189782 202836
rect 237374 202824 237380 202836
rect 189776 202796 237380 202824
rect 189776 202784 189782 202796
rect 237374 202784 237380 202796
rect 237432 202784 237438 202836
rect 2774 201560 2780 201612
rect 2832 201600 2838 201612
rect 4890 201600 4896 201612
rect 2832 201572 4896 201600
rect 2832 201560 2838 201572
rect 4890 201560 4896 201572
rect 4948 201560 4954 201612
rect 187970 201492 187976 201544
rect 188028 201532 188034 201544
rect 237374 201532 237380 201544
rect 188028 201504 237380 201532
rect 188028 201492 188034 201504
rect 237374 201492 237380 201504
rect 237432 201492 237438 201544
rect 189902 200064 189908 200116
rect 189960 200104 189966 200116
rect 237374 200104 237380 200116
rect 189960 200076 237380 200104
rect 189960 200064 189966 200076
rect 237374 200064 237380 200076
rect 237432 200064 237438 200116
rect 136542 199520 136548 199572
rect 136600 199560 136606 199572
rect 237466 199560 237472 199572
rect 136600 199532 237472 199560
rect 136600 199520 136606 199532
rect 237466 199520 237472 199532
rect 237524 199520 237530 199572
rect 105998 199452 106004 199504
rect 106056 199492 106062 199504
rect 238294 199492 238300 199504
rect 106056 199464 238300 199492
rect 106056 199452 106062 199464
rect 238294 199452 238300 199464
rect 238352 199452 238358 199504
rect 103698 199384 103704 199436
rect 103756 199424 103762 199436
rect 188522 199424 188528 199436
rect 103756 199396 188528 199424
rect 103756 199384 103762 199396
rect 188522 199384 188528 199396
rect 188580 199384 188586 199436
rect 150986 199316 150992 199368
rect 151044 199356 151050 199368
rect 235626 199356 235632 199368
rect 151044 199328 235632 199356
rect 151044 199316 151050 199328
rect 235626 199316 235632 199328
rect 235684 199316 235690 199368
rect 86218 199248 86224 199300
rect 86276 199288 86282 199300
rect 187970 199288 187976 199300
rect 86276 199260 187976 199288
rect 86276 199248 86282 199260
rect 187970 199248 187976 199260
rect 188028 199248 188034 199300
rect 83458 199180 83464 199232
rect 83516 199220 83522 199232
rect 187050 199220 187056 199232
rect 83516 199192 187056 199220
rect 83516 199180 83522 199192
rect 187050 199180 187056 199192
rect 187108 199180 187114 199232
rect 82538 199112 82544 199164
rect 82596 199152 82602 199164
rect 187234 199152 187240 199164
rect 82596 199124 187240 199152
rect 82596 199112 82602 199124
rect 187234 199112 187240 199124
rect 187292 199112 187298 199164
rect 81342 199044 81348 199096
rect 81400 199084 81406 199096
rect 187418 199084 187424 199096
rect 81400 199056 187424 199084
rect 81400 199044 81406 199056
rect 187418 199044 187424 199056
rect 187476 199044 187482 199096
rect 77754 198976 77760 199028
rect 77812 199016 77818 199028
rect 187510 199016 187516 199028
rect 77812 198988 187516 199016
rect 77812 198976 77818 198988
rect 187510 198976 187516 198988
rect 187568 198976 187574 199028
rect 71866 198908 71872 198960
rect 71924 198948 71930 198960
rect 188246 198948 188252 198960
rect 71924 198920 188252 198948
rect 71924 198908 71930 198920
rect 188246 198908 188252 198920
rect 188304 198908 188310 198960
rect 91186 198840 91192 198892
rect 91244 198880 91250 198892
rect 238478 198880 238484 198892
rect 91244 198852 238484 198880
rect 91244 198840 91250 198852
rect 238478 198840 238484 198852
rect 238536 198840 238542 198892
rect 88610 198772 88616 198824
rect 88668 198812 88674 198824
rect 237926 198812 237932 198824
rect 88668 198784 237932 198812
rect 88668 198772 88674 198784
rect 237926 198772 237932 198784
rect 237984 198772 237990 198824
rect 78858 198704 78864 198756
rect 78916 198744 78922 198756
rect 228450 198744 228456 198756
rect 78916 198716 228456 198744
rect 78916 198704 78922 198716
rect 228450 198704 228456 198716
rect 228508 198704 228514 198756
rect 84562 198636 84568 198688
rect 84620 198676 84626 198688
rect 238662 198676 238668 198688
rect 84620 198648 238668 198676
rect 84620 198636 84626 198648
rect 238662 198636 238668 198648
rect 238720 198636 238726 198688
rect 88242 198568 88248 198620
rect 88300 198608 88306 198620
rect 238386 198608 238392 198620
rect 88300 198580 238392 198608
rect 88300 198568 88306 198580
rect 238386 198568 238392 198580
rect 238444 198568 238450 198620
rect 93578 198500 93584 198552
rect 93636 198540 93642 198552
rect 238018 198540 238024 198552
rect 93636 198512 238024 198540
rect 93636 198500 93642 198512
rect 238018 198500 238024 198512
rect 238076 198500 238082 198552
rect 93946 198432 93952 198484
rect 94004 198472 94010 198484
rect 235902 198472 235908 198484
rect 94004 198444 235908 198472
rect 94004 198432 94010 198444
rect 235902 198432 235908 198444
rect 235960 198432 235966 198484
rect 80146 198364 80152 198416
rect 80204 198404 80210 198416
rect 105998 198404 106004 198416
rect 80204 198376 106004 198404
rect 80204 198364 80210 198376
rect 105998 198364 106004 198376
rect 106056 198364 106062 198416
rect 106090 198364 106096 198416
rect 106148 198404 106154 198416
rect 238570 198404 238576 198416
rect 106148 198376 238576 198404
rect 106148 198364 106154 198376
rect 238570 198364 238576 198376
rect 238628 198364 238634 198416
rect 95970 198296 95976 198348
rect 96028 198336 96034 198348
rect 188982 198336 188988 198348
rect 96028 198308 188988 198336
rect 96028 198296 96034 198308
rect 188982 198296 188988 198308
rect 189040 198296 189046 198348
rect 98362 198228 98368 198280
rect 98420 198268 98426 198280
rect 188706 198268 188712 198280
rect 98420 198240 188712 198268
rect 98420 198228 98426 198240
rect 188706 198228 188712 198240
rect 188764 198228 188770 198280
rect 76650 198160 76656 198212
rect 76708 198200 76714 198212
rect 136542 198200 136548 198212
rect 76708 198172 136548 198200
rect 76708 198160 76714 198172
rect 136542 198160 136548 198172
rect 136600 198160 136606 198212
rect 148594 198160 148600 198212
rect 148652 198200 148658 198212
rect 235810 198200 235816 198212
rect 148652 198172 235816 198200
rect 148652 198160 148658 198172
rect 235810 198160 235816 198172
rect 235868 198160 235874 198212
rect 100938 198092 100944 198144
rect 100996 198132 101002 198144
rect 188614 198132 188620 198144
rect 100996 198104 188620 198132
rect 100996 198092 101002 198104
rect 188614 198092 188620 198104
rect 188672 198092 188678 198144
rect 123570 198024 123576 198076
rect 123628 198064 123634 198076
rect 188430 198064 188436 198076
rect 123628 198036 188436 198064
rect 123628 198024 123634 198036
rect 188430 198024 188436 198036
rect 188488 198024 188494 198076
rect 70578 197956 70584 198008
rect 70636 197996 70642 198008
rect 237374 197996 237380 198008
rect 70636 197968 237380 197996
rect 70636 197956 70642 197968
rect 237374 197956 237380 197968
rect 237432 197956 237438 198008
rect 99834 197888 99840 197940
rect 99892 197928 99898 197940
rect 128354 197928 128360 197940
rect 99892 197900 128360 197928
rect 99892 197888 99898 197900
rect 128354 197888 128360 197900
rect 128412 197888 128418 197940
rect 128538 197888 128544 197940
rect 128596 197928 128602 197940
rect 188338 197928 188344 197940
rect 128596 197900 188344 197928
rect 128596 197888 128602 197900
rect 188338 197888 188344 197900
rect 188396 197888 188402 197940
rect 130930 197820 130936 197872
rect 130988 197860 130994 197872
rect 188798 197860 188804 197872
rect 130988 197832 188804 197860
rect 130988 197820 130994 197832
rect 188798 197820 188804 197832
rect 188856 197820 188862 197872
rect 136082 197752 136088 197804
rect 136140 197792 136146 197804
rect 188890 197792 188896 197804
rect 136140 197764 188896 197792
rect 136140 197752 136146 197764
rect 188890 197752 188896 197764
rect 188948 197752 188954 197804
rect 173434 197276 173440 197328
rect 173492 197316 173498 197328
rect 194042 197316 194048 197328
rect 173492 197288 194048 197316
rect 173492 197276 173498 197288
rect 194042 197276 194048 197288
rect 194100 197276 194106 197328
rect 232590 197276 232596 197328
rect 232648 197316 232654 197328
rect 237374 197316 237380 197328
rect 232648 197288 237380 197316
rect 232648 197276 232654 197288
rect 237374 197276 237380 197288
rect 237432 197276 237438 197328
rect 173250 197208 173256 197260
rect 173308 197248 173314 197260
rect 192754 197248 192760 197260
rect 173308 197220 192760 197248
rect 173308 197208 173314 197220
rect 192754 197208 192760 197220
rect 192812 197208 192818 197260
rect 47762 197140 47768 197192
rect 47820 197180 47826 197192
rect 191466 197180 191472 197192
rect 47820 197152 191472 197180
rect 47820 197140 47826 197152
rect 191466 197140 191472 197152
rect 191524 197140 191530 197192
rect 48038 197072 48044 197124
rect 48096 197112 48102 197124
rect 191282 197112 191288 197124
rect 48096 197084 191288 197112
rect 48096 197072 48102 197084
rect 191282 197072 191288 197084
rect 191340 197072 191346 197124
rect 105906 197004 105912 197056
rect 105964 197044 105970 197056
rect 235718 197044 235724 197056
rect 105964 197016 235724 197044
rect 105964 197004 105970 197016
rect 235718 197004 235724 197016
rect 235776 197004 235782 197056
rect 107010 196936 107016 196988
rect 107068 196976 107074 196988
rect 235534 196976 235540 196988
rect 107068 196948 235540 196976
rect 107068 196936 107074 196948
rect 235534 196936 235540 196948
rect 235592 196936 235598 196988
rect 85850 196868 85856 196920
rect 85908 196908 85914 196920
rect 195606 196908 195612 196920
rect 85908 196880 195612 196908
rect 85908 196868 85914 196880
rect 195606 196868 195612 196880
rect 195664 196868 195670 196920
rect 87414 196800 87420 196852
rect 87472 196840 87478 196852
rect 191558 196840 191564 196852
rect 87472 196812 191564 196840
rect 87472 196800 87478 196812
rect 191558 196800 191564 196812
rect 191616 196800 191622 196852
rect 90910 196732 90916 196784
rect 90968 196772 90974 196784
rect 189994 196772 190000 196784
rect 90968 196744 190000 196772
rect 90968 196732 90974 196744
rect 189994 196732 190000 196744
rect 190052 196732 190058 196784
rect 92842 196664 92848 196716
rect 92900 196704 92906 196716
rect 191374 196704 191380 196716
rect 92900 196676 191380 196704
rect 92900 196664 92906 196676
rect 191374 196664 191380 196676
rect 191432 196664 191438 196716
rect 102226 196596 102232 196648
rect 102284 196636 102290 196648
rect 189810 196636 189816 196648
rect 102284 196608 189816 196636
rect 102284 196596 102290 196608
rect 189810 196596 189816 196608
rect 189868 196596 189874 196648
rect 108482 196528 108488 196580
rect 108540 196568 108546 196580
rect 186958 196568 186964 196580
rect 108540 196540 186964 196568
rect 108540 196528 108546 196540
rect 186958 196528 186964 196540
rect 187016 196528 187022 196580
rect 89530 196460 89536 196512
rect 89588 196500 89594 196512
rect 238202 196500 238208 196512
rect 89588 196472 238208 196500
rect 89588 196460 89594 196472
rect 238202 196460 238208 196472
rect 238260 196460 238266 196512
rect 92290 196392 92296 196444
rect 92348 196432 92354 196444
rect 238110 196432 238116 196444
rect 92348 196404 238116 196432
rect 92348 196392 92354 196404
rect 238110 196392 238116 196404
rect 238168 196392 238174 196444
rect 189074 195984 189080 196036
rect 189132 196024 189138 196036
rect 237466 196024 237472 196036
rect 189132 195996 237472 196024
rect 189132 195984 189138 195996
rect 237466 195984 237472 195996
rect 237524 195984 237530 196036
rect 75730 195916 75736 195968
rect 75788 195956 75794 195968
rect 237374 195956 237380 195968
rect 75788 195928 237380 195956
rect 75788 195916 75794 195928
rect 237374 195916 237380 195928
rect 237432 195916 237438 195968
rect 83734 195848 83740 195900
rect 83792 195888 83798 195900
rect 189074 195888 189080 195900
rect 83792 195860 189080 195888
rect 83792 195848 83798 195860
rect 189074 195848 189080 195860
rect 189132 195848 189138 195900
rect 111058 195780 111064 195832
rect 111116 195820 111122 195832
rect 193950 195820 193956 195832
rect 111116 195792 193956 195820
rect 111116 195780 111122 195792
rect 193950 195780 193956 195792
rect 194008 195780 194014 195832
rect 113634 195712 113640 195764
rect 113692 195752 113698 195764
rect 195514 195752 195520 195764
rect 113692 195724 195520 195752
rect 113692 195712 113698 195724
rect 195514 195712 195520 195724
rect 195572 195712 195578 195764
rect 153378 195644 153384 195696
rect 153436 195684 153442 195696
rect 235350 195684 235356 195696
rect 153436 195656 235356 195684
rect 153436 195644 153442 195656
rect 235350 195644 235356 195656
rect 235408 195644 235414 195696
rect 116210 195576 116216 195628
rect 116268 195616 116274 195628
rect 195422 195616 195428 195628
rect 116268 195588 195428 195616
rect 116268 195576 116274 195588
rect 195422 195576 195428 195588
rect 195480 195576 195486 195628
rect 155954 195508 155960 195560
rect 156012 195548 156018 195560
rect 235258 195548 235264 195560
rect 156012 195520 235264 195548
rect 156012 195508 156018 195520
rect 235258 195508 235264 195520
rect 235316 195508 235322 195560
rect 118418 195440 118424 195492
rect 118476 195480 118482 195492
rect 195330 195480 195336 195492
rect 118476 195452 195336 195480
rect 118476 195440 118482 195452
rect 195330 195440 195336 195452
rect 195388 195440 195394 195492
rect 120994 195372 121000 195424
rect 121052 195412 121058 195424
rect 196710 195412 196716 195424
rect 121052 195384 196716 195412
rect 121052 195372 121058 195384
rect 196710 195372 196716 195384
rect 196768 195372 196774 195424
rect 126146 195304 126152 195356
rect 126204 195344 126210 195356
rect 196618 195344 196624 195356
rect 126204 195316 196624 195344
rect 126204 195304 126210 195316
rect 196618 195304 196624 195316
rect 196676 195304 196682 195356
rect 133506 195236 133512 195288
rect 133564 195276 133570 195288
rect 197998 195276 198004 195288
rect 133564 195248 198004 195276
rect 133564 195236 133570 195248
rect 197998 195236 198004 195248
rect 198056 195236 198062 195288
rect 146018 195168 146024 195220
rect 146076 195208 146082 195220
rect 192662 195208 192668 195220
rect 146076 195180 192668 195208
rect 146076 195168 146082 195180
rect 192662 195168 192668 195180
rect 192720 195168 192726 195220
rect 49510 194488 49516 194540
rect 49568 194528 49574 194540
rect 237466 194528 237472 194540
rect 49568 194500 237472 194528
rect 49568 194488 49574 194500
rect 237466 194488 237472 194500
rect 237524 194488 237530 194540
rect 198090 194420 198096 194472
rect 198148 194460 198154 194472
rect 237374 194460 237380 194472
rect 198148 194432 237380 194460
rect 198148 194420 198154 194432
rect 237374 194420 237380 194432
rect 237432 194420 237438 194472
rect 69842 193128 69848 193180
rect 69900 193168 69906 193180
rect 237374 193168 237380 193180
rect 69900 193140 237380 193168
rect 69900 193128 69906 193140
rect 237374 193128 237380 193140
rect 237432 193128 237438 193180
rect 499114 191836 499120 191888
rect 499172 191876 499178 191888
rect 579982 191876 579988 191888
rect 499172 191848 579988 191876
rect 499172 191836 499178 191848
rect 579982 191836 579988 191848
rect 580040 191836 580046 191888
rect 81066 191768 81072 191820
rect 81124 191808 81130 191820
rect 237374 191808 237380 191820
rect 81124 191780 237380 191808
rect 81124 191768 81130 191780
rect 237374 191768 237380 191780
rect 237432 191768 237438 191820
rect 232498 191700 232504 191752
rect 232556 191740 232562 191752
rect 237466 191740 237472 191752
rect 232556 191712 237472 191740
rect 232556 191700 232562 191712
rect 237466 191700 237472 191712
rect 237524 191700 237530 191752
rect 74350 190408 74356 190460
rect 74408 190448 74414 190460
rect 237374 190448 237380 190460
rect 74408 190420 237380 190448
rect 74408 190408 74414 190420
rect 237374 190408 237380 190420
rect 237432 190408 237438 190460
rect 192570 190340 192576 190392
rect 192628 190380 192634 190392
rect 237466 190380 237472 190392
rect 192628 190352 237472 190380
rect 192628 190340 192634 190352
rect 237466 190340 237472 190352
rect 237524 190340 237530 190392
rect 67542 188980 67548 189032
rect 67600 189020 67606 189032
rect 237374 189020 237380 189032
rect 67600 188992 237380 189020
rect 67600 188980 67606 188992
rect 237374 188980 237380 188992
rect 237432 188980 237438 189032
rect 68922 187620 68928 187672
rect 68980 187660 68986 187672
rect 237374 187660 237380 187672
rect 68980 187632 237380 187660
rect 68980 187620 68986 187632
rect 237374 187620 237380 187632
rect 237432 187620 237438 187672
rect 78582 186260 78588 186312
rect 78640 186300 78646 186312
rect 237374 186300 237380 186312
rect 78640 186272 237380 186300
rect 78640 186260 78646 186272
rect 237374 186260 237380 186272
rect 237432 186260 237438 186312
rect 580902 185784 580908 185836
rect 580960 185784 580966 185836
rect 580810 185580 580816 185632
rect 580868 185620 580874 185632
rect 580920 185620 580948 185784
rect 580868 185592 580948 185620
rect 580868 185580 580874 185592
rect 74442 184832 74448 184884
rect 74500 184872 74506 184884
rect 237374 184872 237380 184884
rect 74500 184844 237380 184872
rect 74500 184832 74506 184844
rect 237374 184832 237380 184844
rect 237432 184832 237438 184884
rect 192478 184764 192484 184816
rect 192536 184804 192542 184816
rect 237466 184804 237472 184816
rect 192536 184776 237472 184804
rect 192536 184764 192542 184776
rect 237466 184764 237472 184776
rect 237524 184764 237530 184816
rect 66162 183472 66168 183524
rect 66220 183512 66226 183524
rect 237374 183512 237380 183524
rect 66220 183484 237380 183512
rect 66220 183472 66226 183484
rect 237374 183472 237380 183484
rect 237432 183472 237438 183524
rect 49418 182792 49424 182844
rect 49476 182832 49482 182844
rect 237558 182832 237564 182844
rect 49476 182804 237564 182832
rect 49476 182792 49482 182804
rect 237558 182792 237564 182804
rect 237616 182792 237622 182844
rect 47578 182656 47584 182708
rect 47636 182696 47642 182708
rect 48222 182696 48228 182708
rect 47636 182668 48228 182696
rect 47636 182656 47642 182668
rect 48222 182656 48228 182668
rect 48280 182656 48286 182708
rect 48222 182180 48228 182232
rect 48280 182220 48286 182232
rect 88058 182220 88064 182232
rect 48280 182192 88064 182220
rect 48280 182180 48286 182192
rect 88058 182180 88064 182192
rect 88116 182180 88122 182232
rect 49326 182112 49332 182164
rect 49384 182152 49390 182164
rect 237374 182152 237380 182164
rect 49384 182124 237380 182152
rect 49384 182112 49390 182124
rect 237374 182112 237380 182124
rect 237432 182112 237438 182164
rect 215938 182044 215944 182096
rect 215996 182084 216002 182096
rect 237466 182084 237472 182096
rect 215996 182056 237472 182084
rect 215996 182044 216002 182056
rect 237466 182044 237472 182056
rect 237524 182044 237530 182096
rect 23474 181500 23480 181552
rect 23532 181540 23538 181552
rect 237374 181540 237380 181552
rect 23532 181512 237380 181540
rect 23532 181500 23538 181512
rect 237374 181500 237380 181512
rect 237432 181500 237438 181552
rect 3694 181432 3700 181484
rect 3752 181472 3758 181484
rect 238754 181472 238760 181484
rect 3752 181444 238760 181472
rect 3752 181432 3758 181444
rect 238754 181432 238760 181444
rect 238812 181432 238818 181484
rect 218054 180208 218060 180260
rect 218112 180248 218118 180260
rect 366542 180248 366548 180260
rect 218112 180220 366548 180248
rect 218112 180208 218118 180220
rect 366542 180208 366548 180220
rect 366600 180208 366606 180260
rect 367002 180208 367008 180260
rect 367060 180248 367066 180260
rect 580350 180248 580356 180260
rect 367060 180220 580356 180248
rect 367060 180208 367066 180220
rect 580350 180208 580356 180220
rect 580408 180208 580414 180260
rect 300118 180140 300124 180192
rect 300176 180180 300182 180192
rect 580074 180180 580080 180192
rect 300176 180152 580080 180180
rect 300176 180140 300182 180152
rect 580074 180140 580080 180152
rect 580132 180140 580138 180192
rect 3786 180072 3792 180124
rect 3844 180112 3850 180124
rect 435266 180112 435272 180124
rect 3844 180084 435272 180112
rect 3844 180072 3850 180084
rect 435266 180072 435272 180084
rect 435324 180072 435330 180124
rect 233878 179800 233884 179852
rect 233936 179840 233942 179852
rect 386874 179840 386880 179852
rect 233936 179812 386880 179840
rect 233936 179800 233942 179812
rect 386874 179800 386880 179812
rect 386932 179800 386938 179852
rect 239674 179732 239680 179784
rect 239732 179772 239738 179784
rect 432046 179772 432052 179784
rect 239732 179744 432052 179772
rect 239732 179732 239738 179744
rect 432046 179732 432052 179744
rect 432104 179732 432110 179784
rect 346026 179664 346032 179716
rect 346084 179704 346090 179716
rect 542354 179704 542360 179716
rect 346084 179676 542360 179704
rect 346084 179664 346090 179676
rect 542354 179664 542360 179676
rect 542412 179664 542418 179716
rect 239766 179596 239772 179648
rect 239824 179636 239830 179648
rect 438854 179636 438860 179648
rect 239824 179608 438860 179636
rect 239824 179596 239830 179608
rect 438854 179596 438860 179608
rect 438912 179596 438918 179648
rect 191098 179528 191104 179580
rect 191156 179568 191162 179580
rect 393774 179568 393780 179580
rect 191156 179540 393780 179568
rect 191156 179528 191162 179540
rect 393774 179528 393780 179540
rect 393832 179528 393838 179580
rect 239858 179460 239864 179512
rect 239916 179500 239922 179512
rect 445846 179500 445852 179512
rect 239916 179472 445852 179500
rect 239916 179460 239922 179472
rect 445846 179460 445852 179472
rect 445904 179460 445910 179512
rect 3510 179392 3516 179444
rect 3568 179432 3574 179444
rect 421558 179432 421564 179444
rect 3568 179404 421564 179432
rect 3568 179392 3574 179404
rect 421558 179392 421564 179404
rect 421616 179392 421622 179444
rect 3878 179324 3884 179376
rect 3936 179364 3942 179376
rect 483934 179364 483940 179376
rect 3936 179336 483940 179364
rect 3936 179324 3942 179336
rect 483934 179324 483940 179336
rect 483992 179324 483998 179376
rect 3602 179256 3608 179308
rect 3660 179296 3666 179308
rect 428458 179296 428464 179308
rect 3660 179268 428464 179296
rect 3660 179256 3666 179268
rect 428458 179256 428464 179268
rect 428516 179256 428522 179308
rect 46198 179188 46204 179240
rect 46256 179228 46262 179240
rect 459646 179228 459652 179240
rect 46256 179200 459652 179228
rect 46256 179188 46262 179200
rect 459646 179188 459652 179200
rect 459704 179188 459710 179240
rect 43438 179120 43444 179172
rect 43496 179160 43502 179172
rect 452746 179160 452752 179172
rect 43496 179132 452752 179160
rect 43496 179120 43502 179132
rect 452746 179120 452752 179132
rect 452804 179120 452810 179172
rect 325234 179052 325240 179104
rect 325292 179092 325298 179104
rect 580534 179092 580540 179104
rect 325292 179064 580540 179092
rect 325292 179052 325298 179064
rect 580534 179052 580540 179064
rect 580592 179052 580598 179104
rect 335078 178984 335084 179036
rect 335136 179024 335142 179036
rect 580626 179024 580632 179036
rect 335136 178996 580632 179024
rect 335136 178984 335142 178996
rect 580626 178984 580632 178996
rect 580684 178984 580690 179036
rect 236638 178916 236644 178968
rect 236696 178956 236702 178968
rect 473538 178956 473544 178968
rect 236696 178928 473544 178956
rect 236696 178916 236702 178928
rect 473538 178916 473544 178928
rect 473596 178916 473602 178968
rect 483934 178916 483940 178968
rect 483992 178956 483998 178968
rect 580074 178956 580080 178968
rect 483992 178928 580080 178956
rect 483992 178916 483998 178928
rect 580074 178916 580080 178928
rect 580132 178916 580138 178968
rect 240410 178848 240416 178900
rect 240468 178888 240474 178900
rect 348234 178888 348240 178900
rect 240468 178860 348240 178888
rect 240468 178848 240474 178860
rect 348234 178848 348240 178860
rect 348292 178848 348298 178900
rect 349522 178848 349528 178900
rect 349580 178888 349586 178900
rect 580258 178888 580264 178900
rect 349580 178860 580264 178888
rect 349580 178848 349586 178860
rect 580258 178848 580264 178860
rect 580316 178848 580322 178900
rect 239950 178780 239956 178832
rect 240008 178820 240014 178832
rect 295334 178820 295340 178832
rect 240008 178792 295340 178820
rect 240008 178780 240014 178792
rect 295334 178780 295340 178792
rect 295392 178780 295398 178832
rect 307662 178780 307668 178832
rect 307720 178820 307726 178832
rect 498930 178820 498936 178832
rect 307720 178792 498936 178820
rect 307720 178780 307726 178792
rect 498930 178780 498936 178792
rect 498988 178780 498994 178832
rect 239306 178712 239312 178764
rect 239364 178752 239370 178764
rect 311158 178752 311164 178764
rect 239364 178724 311164 178752
rect 239364 178712 239370 178724
rect 311158 178712 311164 178724
rect 311216 178712 311222 178764
rect 318242 178712 318248 178764
rect 318300 178752 318306 178764
rect 498838 178752 498844 178764
rect 318300 178724 498844 178752
rect 318300 178712 318306 178724
rect 498838 178712 498844 178724
rect 498896 178712 498902 178764
rect 3418 178644 3424 178696
rect 3476 178684 3482 178696
rect 380894 178684 380900 178696
rect 3476 178656 380900 178684
rect 3476 178644 3482 178656
rect 380894 178644 380900 178656
rect 380952 178644 380958 178696
rect 398098 178644 398104 178696
rect 398156 178684 398162 178696
rect 580810 178684 580816 178696
rect 398156 178656 580816 178684
rect 398156 178644 398162 178656
rect 580810 178644 580816 178656
rect 580868 178644 580874 178696
rect 239582 178576 239588 178628
rect 239640 178616 239646 178628
rect 404354 178616 404360 178628
rect 239640 178588 404360 178616
rect 239640 178576 239646 178588
rect 404354 178576 404360 178588
rect 404412 178576 404418 178628
rect 239398 178508 239404 178560
rect 239456 178548 239462 178560
rect 397454 178548 397460 178560
rect 239456 178520 397460 178548
rect 239456 178508 239462 178520
rect 397454 178508 397460 178520
rect 397512 178508 397518 178560
rect 363322 178440 363328 178492
rect 363380 178480 363386 178492
rect 500218 178480 500224 178492
rect 363380 178452 500224 178480
rect 363380 178440 363386 178452
rect 500218 178440 500224 178452
rect 500276 178440 500282 178492
rect 490926 178168 490932 178220
rect 490984 178208 490990 178220
rect 492674 178208 492680 178220
rect 490984 178180 492680 178208
rect 490984 178168 490990 178180
rect 492674 178168 492680 178180
rect 492732 178168 492738 178220
rect 380986 178032 380992 178084
rect 381044 178072 381050 178084
rect 580166 178072 580172 178084
rect 381044 178044 580172 178072
rect 381044 178032 381050 178044
rect 580166 178032 580172 178044
rect 580224 178032 580230 178084
rect 348234 177964 348240 178016
rect 348292 178004 348298 178016
rect 372982 178004 372988 178016
rect 348292 177976 372988 178004
rect 348292 177964 348298 177976
rect 372982 177964 372988 177976
rect 373040 177964 373046 178016
rect 380894 177964 380900 178016
rect 380952 178004 380958 178016
rect 414658 178004 414664 178016
rect 380952 177976 414664 178004
rect 380952 177964 380958 177976
rect 414658 177964 414664 177976
rect 414716 177964 414722 178016
rect 435266 177964 435272 178016
rect 435324 178004 435330 178016
rect 449250 178004 449256 178016
rect 435324 177976 449256 178004
rect 435324 177964 435330 177976
rect 449250 177964 449256 177976
rect 449308 177964 449314 178016
rect 4798 177896 4804 177948
rect 4856 177936 4862 177948
rect 463142 177936 463148 177948
rect 4856 177908 463148 177936
rect 4856 177896 4862 177908
rect 463142 177896 463148 177908
rect 463200 177896 463206 177948
rect 88058 177828 88064 177880
rect 88116 177868 88122 177880
rect 241514 177868 241520 177880
rect 88116 177840 241520 177868
rect 88116 177828 88122 177840
rect 241514 177828 241520 177840
rect 241572 177828 241578 177880
rect 293862 177828 293868 177880
rect 293920 177868 293926 177880
rect 300118 177868 300124 177880
rect 293920 177840 300124 177868
rect 293920 177828 293926 177840
rect 300118 177828 300124 177840
rect 300176 177828 300182 177880
rect 328178 177828 328184 177880
rect 328236 177868 328242 177880
rect 580718 177868 580724 177880
rect 328236 177840 580724 177868
rect 328236 177828 328242 177840
rect 580718 177828 580724 177840
rect 580776 177828 580782 177880
rect 341978 177760 341984 177812
rect 342036 177800 342042 177812
rect 580442 177800 580448 177812
rect 342036 177772 580448 177800
rect 342036 177760 342042 177772
rect 580442 177760 580448 177772
rect 580500 177760 580506 177812
rect 228358 177692 228364 177744
rect 228416 177732 228422 177744
rect 455966 177732 455972 177744
rect 228416 177704 455972 177732
rect 228416 177692 228422 177704
rect 455966 177692 455972 177704
rect 456024 177692 456030 177744
rect 456058 177692 456064 177744
rect 456116 177732 456122 177744
rect 477034 177732 477040 177744
rect 456116 177704 477040 177732
rect 456116 177692 456122 177704
rect 477034 177692 477040 177704
rect 477092 177692 477098 177744
rect 276658 177624 276664 177676
rect 276716 177664 276722 177676
rect 500494 177664 500500 177676
rect 276716 177636 500500 177664
rect 276716 177624 276722 177636
rect 500494 177624 500500 177636
rect 500552 177624 500558 177676
rect 283650 177556 283656 177608
rect 283708 177596 283714 177608
rect 500402 177596 500408 177608
rect 283708 177568 500408 177596
rect 283708 177556 283714 177568
rect 500402 177556 500408 177568
rect 500460 177556 500466 177608
rect 297450 177488 297456 177540
rect 297508 177528 297514 177540
rect 501690 177528 501696 177540
rect 297508 177500 501696 177528
rect 297508 177488 297514 177500
rect 501690 177488 501696 177500
rect 501748 177488 501754 177540
rect 304442 177420 304448 177472
rect 304500 177460 304506 177472
rect 501598 177460 501604 177472
rect 304500 177432 501604 177460
rect 304500 177420 304506 177432
rect 501598 177420 501604 177432
rect 501656 177420 501662 177472
rect 290458 177352 290464 177404
rect 290516 177392 290522 177404
rect 483934 177392 483940 177404
rect 290516 177364 483940 177392
rect 290516 177352 290522 177364
rect 483934 177352 483940 177364
rect 483992 177352 483998 177404
rect 1394 177284 1400 177336
rect 1452 177324 1458 177336
rect 244734 177324 244740 177336
rect 1452 177296 244740 177324
rect 1452 177284 1458 177296
rect 244734 177284 244740 177296
rect 244792 177284 244798 177336
rect 377122 177284 377128 177336
rect 377180 177324 377186 177336
rect 485038 177324 485044 177336
rect 377180 177296 485044 177324
rect 377180 177284 377186 177296
rect 485038 177284 485044 177296
rect 485096 177284 485102 177336
rect 240042 177216 240048 177268
rect 240100 177256 240106 177268
rect 390554 177256 390560 177268
rect 240100 177228 390560 177256
rect 240100 177216 240106 177228
rect 390554 177216 390560 177228
rect 390612 177216 390618 177268
rect 321462 177148 321468 177200
rect 321520 177188 321526 177200
rect 398098 177188 398104 177200
rect 321520 177160 398104 177188
rect 321520 177148 321526 177160
rect 398098 177148 398104 177160
rect 398156 177148 398162 177200
rect 4890 177080 4896 177132
rect 4948 177120 4954 177132
rect 470042 177120 470048 177132
rect 4948 177092 470048 177120
rect 4948 177080 4954 177092
rect 470042 177080 470048 177092
rect 470100 177080 470106 177132
rect 269666 177012 269672 177064
rect 269724 177052 269730 177064
rect 380986 177052 380992 177064
rect 269724 177024 380992 177052
rect 269724 177012 269730 177024
rect 380986 177012 380992 177024
rect 381044 177012 381050 177064
rect 493318 176672 493324 176724
rect 493376 176712 493382 176724
rect 498286 176712 498292 176724
rect 493376 176684 498292 176712
rect 493376 176672 493382 176684
rect 498286 176672 498292 176684
rect 498344 176672 498350 176724
rect 6178 176604 6184 176656
rect 6236 176644 6242 176656
rect 480530 176644 480536 176656
rect 6236 176616 480536 176644
rect 6236 176604 6242 176616
rect 480530 176604 480536 176616
rect 480588 176604 480594 176656
rect 311250 176536 311256 176588
rect 311308 176576 311314 176588
rect 580902 176576 580908 176588
rect 311308 176548 580908 176576
rect 311308 176536 311314 176548
rect 580902 176536 580908 176548
rect 580960 176536 580966 176588
rect 286870 176468 286876 176520
rect 286928 176508 286934 176520
rect 499114 176508 499120 176520
rect 286928 176480 499120 176508
rect 286928 176468 286934 176480
rect 499114 176468 499120 176480
rect 499172 176468 499178 176520
rect 300762 176400 300768 176452
rect 300820 176440 300826 176452
rect 499022 176440 499028 176452
rect 300820 176412 499028 176440
rect 300820 176400 300826 176412
rect 499022 176400 499028 176412
rect 499080 176400 499086 176452
rect 314562 176332 314568 176384
rect 314620 176372 314626 176384
rect 500310 176372 500316 176384
rect 314620 176344 500316 176372
rect 314620 176332 314626 176344
rect 500310 176332 500316 176344
rect 500368 176332 500374 176384
rect 359826 176264 359832 176316
rect 359884 176304 359890 176316
rect 490926 176304 490932 176316
rect 359884 176276 490932 176304
rect 359884 176264 359890 176276
rect 490926 176264 490932 176276
rect 490984 176264 490990 176316
rect 295334 176196 295340 176248
rect 295392 176236 295398 176248
rect 383838 176236 383844 176248
rect 295392 176208 383844 176236
rect 295392 176196 295398 176208
rect 383838 176196 383844 176208
rect 383896 176196 383902 176248
rect 311158 176128 311164 176180
rect 311216 176168 311222 176180
rect 366082 176168 366088 176180
rect 311216 176140 366088 176168
rect 311216 176128 311222 176140
rect 366082 176128 366088 176140
rect 366140 176128 366146 176180
rect 278774 153144 278780 153196
rect 278832 153184 278838 153196
rect 580166 153184 580172 153196
rect 278832 153156 580172 153184
rect 278832 153144 278838 153156
rect 580166 153144 580172 153156
rect 580224 153144 580230 153196
rect 3418 150356 3424 150408
rect 3476 150396 3482 150408
rect 456058 150396 456064 150408
rect 3476 150368 456064 150396
rect 3476 150356 3482 150368
rect 456058 150356 456064 150368
rect 456116 150356 456122 150408
rect 3326 141380 3332 141432
rect 3384 141420 3390 141432
rect 487154 141420 487160 141432
rect 3384 141392 487160 141420
rect 3384 141380 3390 141392
rect 487154 141380 487160 141392
rect 487212 141380 487218 141432
rect 262214 139340 262220 139392
rect 262272 139380 262278 139392
rect 580166 139380 580172 139392
rect 262272 139352 580172 139380
rect 262272 139340 262278 139352
rect 580166 139340 580172 139352
rect 580224 139340 580230 139392
rect 271874 113092 271880 113144
rect 271932 113132 271938 113144
rect 579798 113132 579804 113144
rect 271932 113104 579804 113132
rect 271932 113092 271938 113104
rect 579798 113092 579804 113104
rect 579856 113092 579862 113144
rect 255314 100648 255320 100700
rect 255372 100688 255378 100700
rect 580166 100688 580172 100700
rect 255372 100660 580172 100688
rect 255372 100648 255378 100660
rect 580166 100648 580172 100660
rect 580224 100648 580230 100700
rect 3142 85484 3148 85536
rect 3200 85524 3206 85536
rect 489914 85524 489920 85536
rect 3200 85496 489920 85524
rect 3200 85484 3206 85496
rect 489914 85484 489920 85496
rect 489972 85484 489978 85536
rect 264974 73108 264980 73160
rect 265032 73148 265038 73160
rect 580166 73148 580172 73160
rect 265032 73120 580172 73148
rect 265032 73108 265038 73120
rect 580166 73108 580172 73120
rect 580224 73108 580230 73160
rect 248414 60664 248420 60716
rect 248472 60704 248478 60716
rect 580166 60704 580172 60716
rect 248472 60676 580172 60704
rect 248472 60664 248478 60676
rect 580166 60664 580172 60676
rect 580224 60664 580230 60716
rect 3418 45500 3424 45552
rect 3476 45540 3482 45552
rect 494054 45540 494060 45552
rect 3476 45512 494060 45540
rect 3476 45500 3482 45512
rect 494054 45500 494060 45512
rect 494112 45500 494118 45552
rect 258074 33056 258080 33108
rect 258132 33096 258138 33108
rect 580166 33096 580172 33108
rect 258132 33068 580172 33096
rect 258132 33056 258138 33068
rect 580166 33056 580172 33068
rect 580224 33056 580230 33108
rect 3418 6808 3424 6860
rect 3476 6848 3482 6860
rect 493318 6848 493324 6860
rect 3476 6820 493324 6848
rect 3476 6808 3482 6820
rect 493318 6808 493324 6820
rect 493376 6808 493382 6860
rect 251174 6740 251180 6792
rect 251232 6780 251238 6792
rect 580166 6780 580172 6792
rect 251232 6752 580172 6780
rect 251232 6740 251238 6752
rect 580166 6740 580172 6752
rect 580224 6740 580230 6792
rect 566 3408 572 3460
rect 624 3448 630 3460
rect 47578 3448 47584 3460
rect 624 3420 47584 3448
rect 624 3408 630 3420
rect 47578 3408 47584 3420
rect 47636 3408 47642 3460
<< via1 >>
rect 154120 700476 154172 700528
rect 233884 700476 233936 700528
rect 89168 700408 89220 700460
rect 191104 700408 191156 700460
rect 202788 700408 202840 700460
rect 239404 700408 239456 700460
rect 137836 700340 137888 700392
rect 239588 700340 239640 700392
rect 262220 700340 262272 700392
rect 332508 700340 332560 700392
rect 72976 700272 73028 700324
rect 239496 700272 239548 700324
rect 262128 700272 262180 700324
rect 348792 700272 348844 700324
rect 500224 700272 500276 700324
rect 527180 700272 527232 700324
rect 397460 699660 397512 699712
rect 403624 699660 403676 699712
rect 413652 698096 413704 698148
rect 416044 698096 416096 698148
rect 266360 697552 266412 697604
rect 267648 697552 267700 697604
rect 261944 696940 261996 696992
rect 262220 696940 262272 696992
rect 259460 694084 259512 694136
rect 261944 694084 261996 694136
rect 259552 694016 259604 694068
rect 262128 694016 262180 694068
rect 257344 691364 257396 691416
rect 259552 691364 259604 691416
rect 403624 687148 403676 687200
rect 406384 687148 406436 687200
rect 253204 683136 253256 683188
rect 259368 683136 259420 683188
rect 3424 671032 3476 671084
rect 7564 671032 7616 671084
rect 256056 668584 256108 668636
rect 257344 668584 257396 668636
rect 254584 664912 254636 664964
rect 256056 664912 256108 664964
rect 3424 656888 3476 656940
rect 233976 656888 234028 656940
rect 416044 655460 416096 655512
rect 419448 655460 419500 655512
rect 419448 651312 419500 651364
rect 424324 651312 424376 651364
rect 406384 647164 406436 647216
rect 409144 647164 409196 647216
rect 424324 638188 424376 638240
rect 432604 638188 432656 638240
rect 409144 636828 409196 636880
rect 414020 636828 414072 636880
rect 414020 634040 414072 634092
rect 424140 634040 424192 634092
rect 424140 628532 424192 628584
rect 447784 628532 447836 628584
rect 253296 619556 253348 619608
rect 254584 619556 254636 619608
rect 251824 610444 251876 610496
rect 253296 610444 253348 610496
rect 432604 609220 432656 609272
rect 442264 609220 442316 609272
rect 3516 605820 3568 605872
rect 239680 605820 239732 605872
rect 447784 591948 447836 592000
rect 453304 591948 453356 592000
rect 249064 590588 249116 590640
rect 251824 590656 251876 590708
rect 442264 579572 442316 579624
rect 445668 579572 445720 579624
rect 445668 574200 445720 574252
rect 447784 574200 447836 574252
rect 251824 563048 251876 563100
rect 253204 563048 253256 563100
rect 453304 562300 453356 562352
rect 456064 562300 456116 562352
rect 447784 559716 447836 559768
rect 451280 559716 451332 559768
rect 451280 556792 451332 556844
rect 461676 556792 461728 556844
rect 456064 554684 456116 554736
rect 461584 554684 461636 554736
rect 461676 554684 461728 554736
rect 465724 554684 465776 554736
rect 3608 553392 3660 553444
rect 239772 553392 239824 553444
rect 260104 540200 260156 540252
rect 282920 540200 282972 540252
rect 461584 538840 461636 538892
rect 472624 538840 472676 538892
rect 465724 534692 465776 534744
rect 475476 534692 475528 534744
rect 472624 529864 472676 529916
rect 475384 529864 475436 529916
rect 475476 526668 475528 526720
rect 479524 526668 479576 526720
rect 258724 525784 258776 525836
rect 260104 525784 260156 525836
rect 249432 524424 249484 524476
rect 251824 524424 251876 524476
rect 498844 524424 498896 524476
rect 580172 524424 580224 524476
rect 247684 520276 247736 520328
rect 249432 520276 249484 520328
rect 479524 514020 479576 514072
rect 490564 514020 490616 514072
rect 257344 506676 257396 506728
rect 258724 506676 258776 506728
rect 246304 503616 246356 503668
rect 249064 503616 249116 503668
rect 2872 500964 2924 501016
rect 239864 500964 239916 501016
rect 253940 496816 253992 496868
rect 257344 496816 257396 496868
rect 247776 490560 247828 490612
rect 253940 490560 253992 490612
rect 244924 473968 244976 474020
rect 247776 473968 247828 474020
rect 113824 466012 113876 466064
rect 238024 466012 238076 466064
rect 169760 465944 169812 465996
rect 192484 465944 192536 465996
rect 156144 465876 156196 465928
rect 186780 465876 186832 465928
rect 153384 465808 153436 465860
rect 186688 465808 186740 465860
rect 136088 465740 136140 465792
rect 192668 465740 192720 465792
rect 128728 465672 128780 465724
rect 187148 465672 187200 465724
rect 91192 465604 91244 465656
rect 168380 465604 168432 465656
rect 168472 465604 168524 465656
rect 192576 465604 192628 465656
rect 111064 465536 111116 465588
rect 188436 465536 188488 465588
rect 101680 465468 101732 465520
rect 189724 465468 189776 465520
rect 103704 465400 103756 465452
rect 193864 465400 193916 465452
rect 98552 465332 98604 465384
rect 198096 465332 198148 465384
rect 96160 465264 96212 465316
rect 198004 465264 198056 465316
rect 118608 465196 118660 465248
rect 238208 465196 238260 465248
rect 116216 465128 116268 465180
rect 238116 465128 238168 465180
rect 143632 465060 143684 465112
rect 155868 465060 155920 465112
rect 141056 464992 141108 465044
rect 191288 464992 191340 465044
rect 133512 464924 133564 464976
rect 188712 464924 188764 464976
rect 179420 464856 179472 464908
rect 235264 464856 235316 464908
rect 131120 464788 131172 464840
rect 188620 464788 188672 464840
rect 125968 464720 126020 464772
rect 188528 464720 188580 464772
rect 123576 464652 123628 464704
rect 187056 464652 187108 464704
rect 121000 464584 121052 464636
rect 186964 464584 187016 464636
rect 168380 464516 168432 464568
rect 235356 464516 235408 464568
rect 155868 464448 155920 464500
rect 238392 464448 238444 464500
rect 138480 464380 138532 464432
rect 238300 464380 238352 464432
rect 83464 464312 83516 464364
rect 196624 464312 196676 464364
rect 146024 464244 146076 464296
rect 191472 464244 191524 464296
rect 148508 464176 148560 464228
rect 191380 464176 191432 464228
rect 151084 464108 151136 464160
rect 189908 464108 189960 464160
rect 186688 463020 186740 463072
rect 238484 463020 238536 463072
rect 186780 462952 186832 463004
rect 238576 462952 238628 463004
rect 189080 458192 189132 458244
rect 195336 458192 195388 458244
rect 245016 455336 245068 455388
rect 247684 455336 247736 455388
rect 245108 452548 245160 452600
rect 246304 452548 246356 452600
rect 2964 448536 3016 448588
rect 43444 448536 43496 448588
rect 242532 445816 242584 445868
rect 245016 445816 245068 445868
rect 242900 444456 242952 444508
rect 244924 444456 244976 444508
rect 240232 443368 240284 443420
rect 245108 443368 245160 443420
rect 240140 442416 240192 442468
rect 242532 442416 242584 442468
rect 242072 442280 242124 442332
rect 242900 442280 242952 442332
rect 240048 440852 240100 440904
rect 266360 440852 266412 440904
rect 240416 440240 240468 440292
rect 242072 440240 242124 440292
rect 239956 438880 240008 438932
rect 240140 438880 240192 438932
rect 198188 437520 198240 437572
rect 237472 437520 237524 437572
rect 189816 437452 189868 437504
rect 237380 437452 237432 437504
rect 239312 436568 239364 436620
rect 240232 436568 240284 436620
rect 191196 433372 191248 433424
rect 237380 433372 237432 433424
rect 188804 433304 188856 433356
rect 237472 433304 237524 433356
rect 189908 431876 189960 431928
rect 237380 431876 237432 431928
rect 198280 429156 198332 429208
rect 237380 429156 237432 429208
rect 193956 427796 194008 427848
rect 237380 427796 237432 427848
rect 191380 426368 191432 426420
rect 237380 426368 237432 426420
rect 198372 425076 198424 425128
rect 237380 425076 237432 425128
rect 191380 423648 191432 423700
rect 237380 423648 237432 423700
rect 191472 422220 191524 422272
rect 237380 422220 237432 422272
rect 196808 420928 196860 420980
rect 237380 420928 237432 420980
rect 191472 419500 191524 419552
rect 237380 419500 237432 419552
rect 501604 418140 501656 418192
rect 580172 418140 580224 418192
rect 196900 415488 196952 415540
rect 237472 415488 237524 415540
rect 191564 415420 191616 415472
rect 237380 415420 237432 415472
rect 191288 413924 191340 413976
rect 237380 413924 237432 413976
rect 196992 411272 197044 411324
rect 237380 411272 237432 411324
rect 195612 407124 195664 407176
rect 237380 407124 237432 407176
rect 192668 405628 192720 405680
rect 237380 405628 237432 405680
rect 192852 402976 192904 403028
rect 237380 402976 237432 403028
rect 188712 400120 188764 400172
rect 237380 400120 237432 400172
rect 189080 398828 189132 398880
rect 192668 398828 192720 398880
rect 194048 398828 194100 398880
rect 237380 398828 237432 398880
rect 3332 397468 3384 397520
rect 46204 397468 46256 397520
rect 189080 397468 189132 397520
rect 195428 397468 195480 397520
rect 189264 396040 189316 396092
rect 195520 396040 195572 396092
rect 188620 395972 188672 396024
rect 237380 395972 237432 396024
rect 189080 394680 189132 394732
rect 192760 394680 192812 394732
rect 194140 394680 194192 394732
rect 237380 394680 237432 394732
rect 189264 393320 189316 393372
rect 196716 393320 196768 393372
rect 187148 391892 187200 391944
rect 237380 391892 237432 391944
rect 191288 389240 191340 389292
rect 237472 389240 237524 389292
rect 189908 389172 189960 389224
rect 237380 389172 237432 389224
rect 188528 387744 188580 387796
rect 237380 387744 237432 387796
rect 188160 385024 188212 385076
rect 237380 385024 237432 385076
rect 187056 383596 187108 383648
rect 237380 383596 237432 383648
rect 186688 380876 186740 380928
rect 237380 380876 237432 380928
rect 145932 379448 145984 379500
rect 196808 379448 196860 379500
rect 133512 379380 133564 379432
rect 194048 379380 194100 379432
rect 125968 379312 126020 379364
rect 188160 379312 188212 379364
rect 128544 379244 128596 379296
rect 191288 379244 191340 379296
rect 123484 379176 123536 379228
rect 186688 379176 186740 379228
rect 130936 379108 130988 379160
rect 194140 379108 194192 379160
rect 96436 379040 96488 379092
rect 189908 379040 189960 379092
rect 102232 378972 102284 379024
rect 238392 378972 238444 379024
rect 98736 378904 98788 378956
rect 238576 378904 238628 378956
rect 97632 378836 97684 378888
rect 238668 378836 238720 378888
rect 93952 378768 94004 378820
rect 237380 378768 237432 378820
rect 148508 378700 148560 378752
rect 198372 378700 198424 378752
rect 150992 378632 151044 378684
rect 198280 378632 198332 378684
rect 155960 378564 156012 378616
rect 198188 378564 198240 378616
rect 500316 378156 500368 378208
rect 579804 378156 579856 378208
rect 47952 378088 48004 378140
rect 50344 378088 50396 378140
rect 95332 378088 95384 378140
rect 237472 378088 237524 378140
rect 99840 378020 99892 378072
rect 238484 378020 238536 378072
rect 101312 377952 101364 378004
rect 238300 377952 238352 378004
rect 103336 377884 103388 377936
rect 191564 377884 191616 377936
rect 73160 377816 73212 377868
rect 75184 377816 75236 377868
rect 104440 377816 104492 377868
rect 191472 377816 191524 377868
rect 107568 377748 107620 377800
rect 193956 377748 194008 377800
rect 105912 377680 105964 377732
rect 191380 377680 191432 377732
rect 110236 377612 110288 377664
rect 189816 377612 189868 377664
rect 136088 377544 136140 377596
rect 192852 377544 192904 377596
rect 139032 377476 139084 377528
rect 195612 377476 195664 377528
rect 121000 377408 121052 377460
rect 237380 377408 237432 377460
rect 141608 377340 141660 377392
rect 196992 377340 197044 377392
rect 143448 377272 143500 377324
rect 196900 377272 196952 377324
rect 153384 377204 153436 377256
rect 188804 377204 188856 377256
rect 78312 377000 78364 377052
rect 79324 377000 79376 377052
rect 91744 377000 91796 377052
rect 93124 377000 93176 377052
rect 92848 376660 92900 376712
rect 237380 376660 237432 376712
rect 49332 375980 49384 376032
rect 238300 375980 238352 376032
rect 118608 373940 118660 373992
rect 237380 373940 237432 373992
rect 92296 372512 92348 372564
rect 237380 372512 237432 372564
rect 48228 370472 48280 370524
rect 148324 370472 148376 370524
rect 91008 368432 91060 368484
rect 237472 368432 237524 368484
rect 117228 368364 117280 368416
rect 237380 368364 237432 368416
rect 47860 367752 47912 367804
rect 122104 367752 122156 367804
rect 48044 365644 48096 365696
rect 50436 365644 50488 365696
rect 501696 364352 501748 364404
rect 580172 364352 580224 364404
rect 89536 364284 89588 364336
rect 237472 364284 237524 364336
rect 114468 364216 114520 364268
rect 237380 364216 237432 364268
rect 188436 361496 188488 361548
rect 237380 361496 237432 361548
rect 111708 360136 111760 360188
rect 237380 360136 237432 360188
rect 48136 359456 48188 359508
rect 167644 359456 167696 359508
rect 88156 358708 88208 358760
rect 237380 358708 237432 358760
rect 108948 355988 109000 356040
rect 237380 355988 237432 356040
rect 88248 354628 88300 354680
rect 237380 354628 237432 354680
rect 106188 351840 106240 351892
rect 237380 351840 237432 351892
rect 86776 350480 86828 350532
rect 237380 350480 237432 350532
rect 104808 347692 104860 347744
rect 237472 347692 237524 347744
rect 193864 347624 193916 347676
rect 237380 347624 237432 347676
rect 49424 347012 49476 347064
rect 238024 347012 238076 347064
rect 85488 346332 85540 346384
rect 237380 346332 237432 346384
rect 189724 343544 189776 343596
rect 237380 343544 237432 343596
rect 84016 342184 84068 342236
rect 237472 342184 237524 342236
rect 102048 342116 102100 342168
rect 237380 342116 237432 342168
rect 3884 340144 3936 340196
rect 191196 340144 191248 340196
rect 198096 339396 198148 339448
rect 237380 339396 237432 339448
rect 82728 338036 82780 338088
rect 237472 338036 237524 338088
rect 99288 337968 99340 338020
rect 237380 337968 237432 338020
rect 173716 336676 173768 336728
rect 237380 336676 237432 336728
rect 50436 335248 50488 335300
rect 237380 335248 237432 335300
rect 198004 335180 198056 335232
rect 237472 335180 237524 335232
rect 96528 333888 96580 333940
rect 237380 333888 237432 333940
rect 81164 332528 81216 332580
rect 237380 332528 237432 332580
rect 173808 332460 173860 332512
rect 237472 332460 237524 332512
rect 167644 331168 167696 331220
rect 237380 331168 237432 331220
rect 93768 329740 93820 329792
rect 237380 329740 237432 329792
rect 81256 328380 81308 328432
rect 237380 328380 237432 328432
rect 196716 328312 196768 328364
rect 237472 328312 237524 328364
rect 50344 327020 50396 327072
rect 237380 327020 237432 327072
rect 93124 325592 93176 325644
rect 237380 325592 237432 325644
rect 235356 325524 235408 325576
rect 237472 325524 237524 325576
rect 499028 324300 499080 324352
rect 579988 324300 580040 324352
rect 79968 324232 80020 324284
rect 237380 324232 237432 324284
rect 192760 322872 192812 322924
rect 237380 322872 237432 322924
rect 235264 321512 235316 321564
rect 237380 321512 237432 321564
rect 78496 320084 78548 320136
rect 237472 320084 237524 320136
rect 89628 320016 89680 320068
rect 237380 320016 237432 320068
rect 195520 318724 195572 318776
rect 237380 318724 237432 318776
rect 73068 317364 73120 317416
rect 237380 317364 237432 317416
rect 86868 315936 86920 315988
rect 237380 315936 237432 315988
rect 77208 314576 77260 314628
rect 237380 314576 237432 314628
rect 49240 313216 49292 313268
rect 237472 313216 237524 313268
rect 195428 313148 195480 313200
rect 237380 313148 237432 313200
rect 71688 311788 71740 311840
rect 237380 311788 237432 311840
rect 84108 310428 84160 310480
rect 237472 310428 237524 310480
rect 196624 310360 196676 310412
rect 237380 310360 237432 310412
rect 75828 309068 75880 309120
rect 237380 309068 237432 309120
rect 192668 309000 192720 309052
rect 237472 309000 237524 309052
rect 49608 307708 49660 307760
rect 237380 307708 237432 307760
rect 70308 306280 70360 306332
rect 237380 306280 237432 306332
rect 188344 306212 188396 306264
rect 237472 306212 237524 306264
rect 3148 304988 3200 305040
rect 228364 304988 228416 305040
rect 81348 304920 81400 304972
rect 237380 304920 237432 304972
rect 74356 303560 74408 303612
rect 237380 303560 237432 303612
rect 192576 303492 192628 303544
rect 237472 303492 237524 303544
rect 67548 302132 67600 302184
rect 237380 302132 237432 302184
rect 68928 300772 68980 300824
rect 237380 300772 237432 300824
rect 195244 300704 195296 300756
rect 237472 300704 237524 300756
rect 75184 299412 75236 299464
rect 237472 299412 237524 299464
rect 79324 299344 79376 299396
rect 237380 299344 237432 299396
rect 192484 298052 192536 298104
rect 237380 298052 237432 298104
rect 66168 296624 66220 296676
rect 237380 296624 237432 296676
rect 148324 296556 148376 296608
rect 237472 296556 237524 296608
rect 195336 295264 195388 295316
rect 237380 295264 237432 295316
rect 122104 293904 122156 293956
rect 237380 293904 237432 293956
rect 157248 292612 157300 292664
rect 237380 292612 237432 292664
rect 3332 292544 3384 292596
rect 236644 292544 236696 292596
rect 235264 291184 235316 291236
rect 237380 291184 237432 291236
rect 154488 289824 154540 289876
rect 237380 289824 237432 289876
rect 235356 288464 235408 288516
rect 237472 288464 237524 288516
rect 235448 288396 235500 288448
rect 237380 288396 237432 288448
rect 151728 287036 151780 287088
rect 237380 287036 237432 287088
rect 170680 286560 170732 286612
rect 192484 286560 192536 286612
rect 169668 286492 169720 286544
rect 192576 286492 192628 286544
rect 144828 286424 144880 286476
rect 186780 286424 186832 286476
rect 141884 286356 141936 286408
rect 187332 286356 187384 286408
rect 139308 286288 139360 286340
rect 187240 286288 187292 286340
rect 136548 286220 136600 286272
rect 187148 286220 187200 286272
rect 126888 286152 126940 286204
rect 187056 286152 187108 286204
rect 124128 286084 124180 286136
rect 186964 286084 187016 286136
rect 108948 286016 109000 286068
rect 194048 286016 194100 286068
rect 106188 285948 106240 286000
rect 191472 285948 191524 286000
rect 104808 285880 104860 285932
rect 192760 285880 192812 285932
rect 118608 285812 118660 285864
rect 238116 285880 238168 285932
rect 114468 285744 114520 285796
rect 238208 285812 238260 285864
rect 235540 285744 235592 285796
rect 237472 285744 237524 285796
rect 83740 285676 83792 285728
rect 232596 285676 232648 285728
rect 235632 285676 235684 285728
rect 237380 285676 237432 285728
rect 92388 285608 92440 285660
rect 191288 285608 191340 285660
rect 93676 285540 93728 285592
rect 195244 285540 195296 285592
rect 96528 285472 96580 285524
rect 198096 285472 198148 285524
rect 86868 285404 86920 285456
rect 189724 285404 189776 285456
rect 133788 285336 133840 285388
rect 237840 285336 237892 285388
rect 89628 285268 89680 285320
rect 193864 285268 193916 285320
rect 131120 285200 131172 285252
rect 238484 285200 238536 285252
rect 128728 285132 128780 285184
rect 238668 285132 238720 285184
rect 116216 285064 116268 285116
rect 238576 285064 238628 285116
rect 111064 284996 111116 285048
rect 238392 284996 238444 285048
rect 98552 284928 98604 284980
rect 238024 284928 238076 284980
rect 148600 284860 148652 284912
rect 237380 284860 237432 284912
rect 101312 284792 101364 284844
rect 189908 284792 189960 284844
rect 146024 284724 146076 284776
rect 186688 284724 186740 284776
rect 235816 282956 235868 283008
rect 237380 282956 237432 283008
rect 235724 282888 235776 282940
rect 237472 282888 237524 282940
rect 186688 282820 186740 282872
rect 237380 282820 237432 282872
rect 192668 280236 192720 280288
rect 237380 280236 237432 280288
rect 187608 280168 187660 280220
rect 237472 280168 237524 280220
rect 186780 280100 186832 280152
rect 237380 280100 237432 280152
rect 190000 278740 190052 278792
rect 215944 278740 215996 278792
rect 187332 277312 187384 277364
rect 237380 277312 237432 277364
rect 189816 274660 189868 274712
rect 237472 274660 237524 274712
rect 187240 274592 187292 274644
rect 237380 274592 237432 274644
rect 499028 271872 499080 271924
rect 579804 271872 579856 271924
rect 187148 271804 187200 271856
rect 237380 271804 237432 271856
rect 198004 267724 198056 267776
rect 237380 267724 237432 267776
rect 188344 262216 188396 262268
rect 237380 262216 237432 262268
rect 187056 262148 187108 262200
rect 237472 262148 237524 262200
rect 187148 260856 187200 260908
rect 237380 260856 237432 260908
rect 196624 259496 196676 259548
rect 237380 259496 237432 259548
rect 187332 259428 187384 259480
rect 237472 259428 237524 259480
rect 186964 259360 187016 259412
rect 237380 259360 237432 259412
rect 500408 258068 500460 258120
rect 579988 258068 580040 258120
rect 235908 256776 235960 256828
rect 237472 256776 237524 256828
rect 188436 256708 188488 256760
rect 237380 256708 237432 256760
rect 2780 254056 2832 254108
rect 4804 254056 4856 254108
rect 196716 253988 196768 254040
rect 237472 253988 237524 254040
rect 191380 253920 191432 253972
rect 237380 253920 237432 253972
rect 195336 251200 195388 251252
rect 237380 251200 237432 251252
rect 195428 249772 195480 249824
rect 237380 249772 237432 249824
rect 190000 248412 190052 248464
rect 237380 248412 237432 248464
rect 195520 247052 195572 247104
rect 237380 247052 237432 247104
rect 193956 244264 194008 244316
rect 237380 244264 237432 244316
rect 194048 242836 194100 242888
rect 237380 242836 237432 242888
rect 186964 241476 187016 241528
rect 237380 241476 237432 241528
rect 3148 240320 3200 240372
rect 6184 240320 6236 240372
rect 191564 240116 191616 240168
rect 237380 240116 237432 240168
rect 191472 238688 191524 238740
rect 237380 238688 237432 238740
rect 195612 235968 195664 236020
rect 237380 235968 237432 236020
rect 192760 234540 192812 234592
rect 237380 234540 237432 234592
rect 188528 231820 188580 231872
rect 237380 231820 237432 231872
rect 189908 230392 189960 230444
rect 237380 230392 237432 230444
rect 188620 227808 188672 227860
rect 237472 227808 237524 227860
rect 187056 227740 187108 227792
rect 237380 227740 237432 227792
rect 188712 223592 188764 223644
rect 237380 223592 237432 223644
rect 194048 222232 194100 222284
rect 237380 222232 237432 222284
rect 187240 222164 187292 222216
rect 237472 222164 237524 222216
rect 198096 222096 198148 222148
rect 237380 222096 237432 222148
rect 188896 221484 188948 221536
rect 238300 221484 238352 221536
rect 188804 221416 188856 221468
rect 238484 221416 238536 221468
rect 235172 220804 235224 220856
rect 237472 220804 237524 220856
rect 188988 219444 189040 219496
rect 237380 219444 237432 219496
rect 189080 218152 189132 218204
rect 198096 218152 198148 218204
rect 192760 218084 192812 218136
rect 237380 218084 237432 218136
rect 187424 218016 187476 218068
rect 237472 218016 237524 218068
rect 500500 218016 500552 218068
rect 579804 218016 579856 218068
rect 195244 216588 195296 216640
rect 237380 216588 237432 216640
rect 189080 215296 189132 215348
rect 191472 215296 191524 215348
rect 190092 213936 190144 213988
rect 191656 213936 191708 213988
rect 190276 213188 190328 213240
rect 237380 213188 237432 213240
rect 234988 212508 235040 212560
rect 237472 212508 237524 212560
rect 191288 212440 191340 212492
rect 237380 212440 237432 212492
rect 228456 209788 228508 209840
rect 237472 209788 237524 209840
rect 191656 209720 191708 209772
rect 237380 209720 237432 209772
rect 191288 208360 191340 208412
rect 237380 208360 237432 208412
rect 193864 208292 193916 208344
rect 237472 208292 237524 208344
rect 47584 207680 47636 207732
rect 48228 207680 48280 207732
rect 49608 207680 49660 207732
rect 187516 205640 187568 205692
rect 237472 205640 237524 205692
rect 191472 205572 191524 205624
rect 237380 205572 237432 205624
rect 191472 202920 191524 202972
rect 237380 202920 237432 202972
rect 188252 202852 188304 202904
rect 237472 202852 237524 202904
rect 189724 202784 189776 202836
rect 237380 202784 237432 202836
rect 2780 201560 2832 201612
rect 4896 201560 4948 201612
rect 187976 201492 188028 201544
rect 237380 201492 237432 201544
rect 189908 200064 189960 200116
rect 237380 200064 237432 200116
rect 136548 199520 136600 199572
rect 237472 199520 237524 199572
rect 106004 199452 106056 199504
rect 238300 199452 238352 199504
rect 103704 199384 103756 199436
rect 188528 199384 188580 199436
rect 150992 199316 151044 199368
rect 235632 199316 235684 199368
rect 86224 199248 86276 199300
rect 187976 199248 188028 199300
rect 83464 199180 83516 199232
rect 187056 199180 187108 199232
rect 82544 199112 82596 199164
rect 187240 199112 187292 199164
rect 81348 199044 81400 199096
rect 187424 199044 187476 199096
rect 77760 198976 77812 199028
rect 187516 198976 187568 199028
rect 71872 198908 71924 198960
rect 188252 198908 188304 198960
rect 91192 198840 91244 198892
rect 238484 198840 238536 198892
rect 88616 198772 88668 198824
rect 237932 198772 237984 198824
rect 78864 198704 78916 198756
rect 228456 198704 228508 198756
rect 84568 198636 84620 198688
rect 238668 198636 238720 198688
rect 88248 198568 88300 198620
rect 238392 198568 238444 198620
rect 93584 198500 93636 198552
rect 238024 198500 238076 198552
rect 93952 198432 94004 198484
rect 235908 198432 235960 198484
rect 80152 198364 80204 198416
rect 106004 198364 106056 198416
rect 106096 198364 106148 198416
rect 238576 198364 238628 198416
rect 95976 198296 96028 198348
rect 188988 198296 189040 198348
rect 98368 198228 98420 198280
rect 188712 198228 188764 198280
rect 76656 198160 76708 198212
rect 136548 198160 136600 198212
rect 148600 198160 148652 198212
rect 235816 198160 235868 198212
rect 100944 198092 100996 198144
rect 188620 198092 188672 198144
rect 123576 198024 123628 198076
rect 188436 198024 188488 198076
rect 70584 197956 70636 198008
rect 237380 197956 237432 198008
rect 99840 197888 99892 197940
rect 128360 197888 128412 197940
rect 128544 197888 128596 197940
rect 188344 197888 188396 197940
rect 130936 197820 130988 197872
rect 188804 197820 188856 197872
rect 136088 197752 136140 197804
rect 188896 197752 188948 197804
rect 173440 197276 173492 197328
rect 194048 197276 194100 197328
rect 232596 197276 232648 197328
rect 237380 197276 237432 197328
rect 173256 197208 173308 197260
rect 192760 197208 192812 197260
rect 47768 197140 47820 197192
rect 191472 197140 191524 197192
rect 48044 197072 48096 197124
rect 191288 197072 191340 197124
rect 105912 197004 105964 197056
rect 235724 197004 235776 197056
rect 107016 196936 107068 196988
rect 235540 196936 235592 196988
rect 85856 196868 85908 196920
rect 195612 196868 195664 196920
rect 87420 196800 87472 196852
rect 191564 196800 191616 196852
rect 90916 196732 90968 196784
rect 190000 196732 190052 196784
rect 92848 196664 92900 196716
rect 191380 196664 191432 196716
rect 102232 196596 102284 196648
rect 189816 196596 189868 196648
rect 108488 196528 108540 196580
rect 186964 196528 187016 196580
rect 89536 196460 89588 196512
rect 238208 196460 238260 196512
rect 92296 196392 92348 196444
rect 238116 196392 238168 196444
rect 189080 195984 189132 196036
rect 237472 195984 237524 196036
rect 75736 195916 75788 195968
rect 237380 195916 237432 195968
rect 83740 195848 83792 195900
rect 189080 195848 189132 195900
rect 111064 195780 111116 195832
rect 193956 195780 194008 195832
rect 113640 195712 113692 195764
rect 195520 195712 195572 195764
rect 153384 195644 153436 195696
rect 235356 195644 235408 195696
rect 116216 195576 116268 195628
rect 195428 195576 195480 195628
rect 155960 195508 156012 195560
rect 235264 195508 235316 195560
rect 118424 195440 118476 195492
rect 195336 195440 195388 195492
rect 121000 195372 121052 195424
rect 196716 195372 196768 195424
rect 126152 195304 126204 195356
rect 196624 195304 196676 195356
rect 133512 195236 133564 195288
rect 198004 195236 198056 195288
rect 146024 195168 146076 195220
rect 192668 195168 192720 195220
rect 49516 194488 49568 194540
rect 237472 194488 237524 194540
rect 198096 194420 198148 194472
rect 237380 194420 237432 194472
rect 69848 193128 69900 193180
rect 237380 193128 237432 193180
rect 499120 191836 499172 191888
rect 579988 191836 580040 191888
rect 81072 191768 81124 191820
rect 237380 191768 237432 191820
rect 232504 191700 232556 191752
rect 237472 191700 237524 191752
rect 74356 190408 74408 190460
rect 237380 190408 237432 190460
rect 192576 190340 192628 190392
rect 237472 190340 237524 190392
rect 67548 188980 67600 189032
rect 237380 188980 237432 189032
rect 68928 187620 68980 187672
rect 237380 187620 237432 187672
rect 78588 186260 78640 186312
rect 237380 186260 237432 186312
rect 580908 185784 580960 185836
rect 580816 185580 580868 185632
rect 74448 184832 74500 184884
rect 237380 184832 237432 184884
rect 192484 184764 192536 184816
rect 237472 184764 237524 184816
rect 66168 183472 66220 183524
rect 237380 183472 237432 183524
rect 49424 182792 49476 182844
rect 237564 182792 237616 182844
rect 47584 182656 47636 182708
rect 48228 182656 48280 182708
rect 48228 182180 48280 182232
rect 88064 182180 88116 182232
rect 49332 182112 49384 182164
rect 237380 182112 237432 182164
rect 215944 182044 215996 182096
rect 237472 182044 237524 182096
rect 23480 181500 23532 181552
rect 237380 181500 237432 181552
rect 3700 181432 3752 181484
rect 238760 181432 238812 181484
rect 218060 180208 218112 180260
rect 366548 180208 366600 180260
rect 367008 180208 367060 180260
rect 580356 180208 580408 180260
rect 300124 180140 300176 180192
rect 580080 180140 580132 180192
rect 3792 180072 3844 180124
rect 435272 180072 435324 180124
rect 233884 179800 233936 179852
rect 386880 179800 386932 179852
rect 239680 179732 239732 179784
rect 432052 179732 432104 179784
rect 346032 179664 346084 179716
rect 542360 179664 542412 179716
rect 239772 179596 239824 179648
rect 438860 179596 438912 179648
rect 191104 179528 191156 179580
rect 393780 179528 393832 179580
rect 239864 179460 239916 179512
rect 445852 179460 445904 179512
rect 3516 179392 3568 179444
rect 421564 179392 421616 179444
rect 3884 179324 3936 179376
rect 483940 179324 483992 179376
rect 3608 179256 3660 179308
rect 428464 179256 428516 179308
rect 46204 179188 46256 179240
rect 459652 179188 459704 179240
rect 43444 179120 43496 179172
rect 452752 179120 452804 179172
rect 325240 179052 325292 179104
rect 580540 179052 580592 179104
rect 335084 178984 335136 179036
rect 580632 178984 580684 179036
rect 236644 178916 236696 178968
rect 473544 178916 473596 178968
rect 483940 178916 483992 178968
rect 580080 178916 580132 178968
rect 240416 178848 240468 178900
rect 348240 178848 348292 178900
rect 349528 178848 349580 178900
rect 580264 178848 580316 178900
rect 239956 178780 240008 178832
rect 295340 178780 295392 178832
rect 307668 178780 307720 178832
rect 498936 178780 498988 178832
rect 239312 178712 239364 178764
rect 311164 178712 311216 178764
rect 318248 178712 318300 178764
rect 498844 178712 498896 178764
rect 3424 178644 3476 178696
rect 380900 178644 380952 178696
rect 398104 178644 398156 178696
rect 580816 178644 580868 178696
rect 239588 178576 239640 178628
rect 404360 178576 404412 178628
rect 239404 178508 239456 178560
rect 397460 178508 397512 178560
rect 363328 178440 363380 178492
rect 500224 178440 500276 178492
rect 490932 178168 490984 178220
rect 492680 178168 492732 178220
rect 380992 178032 381044 178084
rect 580172 178032 580224 178084
rect 348240 177964 348292 178016
rect 372988 177964 373040 178016
rect 380900 177964 380952 178016
rect 414664 177964 414716 178016
rect 435272 177964 435324 178016
rect 449256 177964 449308 178016
rect 4804 177896 4856 177948
rect 463148 177896 463200 177948
rect 88064 177828 88116 177880
rect 241520 177828 241572 177880
rect 293868 177828 293920 177880
rect 300124 177828 300176 177880
rect 328184 177828 328236 177880
rect 580724 177828 580776 177880
rect 341984 177760 342036 177812
rect 580448 177760 580500 177812
rect 228364 177692 228416 177744
rect 455972 177692 456024 177744
rect 456064 177692 456116 177744
rect 477040 177692 477092 177744
rect 276664 177624 276716 177676
rect 500500 177624 500552 177676
rect 283656 177556 283708 177608
rect 500408 177556 500460 177608
rect 297456 177488 297508 177540
rect 501696 177488 501748 177540
rect 304448 177420 304500 177472
rect 501604 177420 501656 177472
rect 290464 177352 290516 177404
rect 483940 177352 483992 177404
rect 1400 177284 1452 177336
rect 244740 177284 244792 177336
rect 377128 177284 377180 177336
rect 485044 177284 485096 177336
rect 240048 177216 240100 177268
rect 390560 177216 390612 177268
rect 321468 177148 321520 177200
rect 398104 177148 398156 177200
rect 4896 177080 4948 177132
rect 470048 177080 470100 177132
rect 269672 177012 269724 177064
rect 380992 177012 381044 177064
rect 493324 176672 493376 176724
rect 498292 176672 498344 176724
rect 6184 176604 6236 176656
rect 480536 176604 480588 176656
rect 311256 176536 311308 176588
rect 580908 176536 580960 176588
rect 286876 176468 286928 176520
rect 499120 176468 499172 176520
rect 300768 176400 300820 176452
rect 499028 176400 499080 176452
rect 314568 176332 314620 176384
rect 500316 176332 500368 176384
rect 359832 176264 359884 176316
rect 490932 176264 490984 176316
rect 295340 176196 295392 176248
rect 383844 176196 383896 176248
rect 311164 176128 311216 176180
rect 366088 176128 366140 176180
rect 278780 153144 278832 153196
rect 580172 153144 580224 153196
rect 3424 150356 3476 150408
rect 456064 150356 456116 150408
rect 3332 141380 3384 141432
rect 487160 141380 487212 141432
rect 262220 139340 262272 139392
rect 580172 139340 580224 139392
rect 271880 113092 271932 113144
rect 579804 113092 579856 113144
rect 255320 100648 255372 100700
rect 580172 100648 580224 100700
rect 3148 85484 3200 85536
rect 489920 85484 489972 85536
rect 264980 73108 265032 73160
rect 580172 73108 580224 73160
rect 248420 60664 248472 60716
rect 580172 60664 580224 60716
rect 3424 45500 3476 45552
rect 494060 45500 494112 45552
rect 258080 33056 258132 33108
rect 580172 33056 580224 33108
rect 3424 6808 3476 6860
rect 493324 6808 493376 6860
rect 251180 6740 251232 6792
rect 580172 6740 580224 6792
rect 572 3408 624 3460
rect 47584 3408 47636 3460
<< metal2 >>
rect 8086 703520 8198 704960
rect 23492 703582 24164 703610
rect 8128 700369 8156 703520
rect 8114 700360 8170 700369
rect 8114 700295 8170 700304
rect 3422 671256 3478 671265
rect 3422 671191 3478 671200
rect 3436 671090 3464 671191
rect 3424 671084 3476 671090
rect 3424 671026 3476 671032
rect 7564 671084 7616 671090
rect 7564 671026 7616 671032
rect 3422 658200 3478 658209
rect 3422 658135 3478 658144
rect 3436 656946 3464 658135
rect 3424 656940 3476 656946
rect 3424 656882 3476 656888
rect 3422 619168 3478 619177
rect 3422 619103 3478 619112
rect 2870 501800 2926 501809
rect 2870 501735 2926 501744
rect 2884 501022 2912 501735
rect 2872 501016 2924 501022
rect 2872 500958 2924 500964
rect 2962 449576 3018 449585
rect 2962 449511 3018 449520
rect 2976 448594 3004 449511
rect 2964 448588 3016 448594
rect 2964 448530 3016 448536
rect 3332 397520 3384 397526
rect 3330 397488 3332 397497
rect 3384 397488 3386 397497
rect 3330 397423 3386 397432
rect 3146 306232 3202 306241
rect 3146 306167 3202 306176
rect 3160 305046 3188 306167
rect 3148 305040 3200 305046
rect 3148 304982 3200 304988
rect 3330 293176 3386 293185
rect 3330 293111 3386 293120
rect 3344 292602 3372 293111
rect 3332 292596 3384 292602
rect 3332 292538 3384 292544
rect 2778 254144 2834 254153
rect 2778 254079 2780 254088
rect 2832 254079 2834 254088
rect 2780 254050 2832 254056
rect 3146 241088 3202 241097
rect 3146 241023 3202 241032
rect 3160 240378 3188 241023
rect 3148 240372 3200 240378
rect 3148 240314 3200 240320
rect 2778 201920 2834 201929
rect 2778 201855 2834 201864
rect 2792 201618 2820 201855
rect 2780 201612 2832 201618
rect 2780 201554 2832 201560
rect 3436 178702 3464 619103
rect 3514 606112 3570 606121
rect 3514 606047 3570 606056
rect 3528 605878 3556 606047
rect 3516 605872 3568 605878
rect 3516 605814 3568 605820
rect 3514 566944 3570 566953
rect 3514 566879 3570 566888
rect 3528 179450 3556 566879
rect 3606 553888 3662 553897
rect 3606 553823 3662 553832
rect 3620 553450 3648 553823
rect 3608 553444 3660 553450
rect 3608 553386 3660 553392
rect 3606 514856 3662 514865
rect 3606 514791 3662 514800
rect 3516 179444 3568 179450
rect 3516 179386 3568 179392
rect 3620 179314 3648 514791
rect 3698 462632 3754 462641
rect 3698 462567 3754 462576
rect 3712 181490 3740 462567
rect 3882 410544 3938 410553
rect 3882 410479 3938 410488
rect 3790 358456 3846 358465
rect 3790 358391 3846 358400
rect 3700 181484 3752 181490
rect 3700 181426 3752 181432
rect 3804 180130 3832 358391
rect 3896 340202 3924 410479
rect 3884 340196 3936 340202
rect 3884 340138 3936 340144
rect 4804 254108 4856 254114
rect 4804 254050 4856 254056
rect 3882 188864 3938 188873
rect 3882 188799 3938 188808
rect 3792 180124 3844 180130
rect 3792 180066 3844 180072
rect 3896 179382 3924 188799
rect 3884 179376 3936 179382
rect 3884 179318 3936 179324
rect 3608 179308 3660 179314
rect 3608 179250 3660 179256
rect 3424 178696 3476 178702
rect 3424 178638 3476 178644
rect 4816 177954 4844 254050
rect 6184 240372 6236 240378
rect 6184 240314 6236 240320
rect 4896 201612 4948 201618
rect 4896 201554 4948 201560
rect 4804 177948 4856 177954
rect 4804 177890 4856 177896
rect 1400 177336 1452 177342
rect 1400 177278 1452 177284
rect 572 3460 624 3466
rect 572 3402 624 3408
rect 584 480 612 3402
rect 542 -960 654 480
rect 1412 354 1440 177278
rect 4908 177138 4936 201554
rect 4896 177132 4948 177138
rect 4896 177074 4948 177080
rect 6196 176662 6224 240314
rect 7576 179489 7604 671026
rect 23492 181558 23520 703582
rect 24136 703474 24164 703582
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218072 703582 218836 703610
rect 24320 703474 24348 703520
rect 24136 703446 24348 703474
rect 72988 700330 73016 703520
rect 89180 700466 89208 703520
rect 89168 700460 89220 700466
rect 89168 700402 89220 700408
rect 137848 700398 137876 703520
rect 154132 700534 154160 703520
rect 154120 700528 154172 700534
rect 154120 700470 154172 700476
rect 202800 700466 202828 703520
rect 191104 700460 191156 700466
rect 191104 700402 191156 700408
rect 202788 700460 202840 700466
rect 202788 700402 202840 700408
rect 137836 700392 137888 700398
rect 137836 700334 137888 700340
rect 72976 700324 73028 700330
rect 72976 700266 73028 700272
rect 113824 466064 113876 466070
rect 113824 466006 113876 466012
rect 179418 466032 179474 466041
rect 91192 465656 91244 465662
rect 91192 465598 91244 465604
rect 91204 465225 91232 465598
rect 111064 465588 111116 465594
rect 111064 465530 111116 465536
rect 101680 465520 101732 465526
rect 101680 465462 101732 465468
rect 98552 465384 98604 465390
rect 98552 465326 98604 465332
rect 96160 465316 96212 465322
rect 96160 465258 96212 465264
rect 96172 465225 96200 465258
rect 98564 465225 98592 465326
rect 101692 465225 101720 465462
rect 103704 465452 103756 465458
rect 103704 465394 103756 465400
rect 103716 465225 103744 465394
rect 111076 465225 111104 465530
rect 113836 465225 113864 466006
rect 169760 465996 169812 466002
rect 179418 465967 179474 465976
rect 169760 465938 169812 465944
rect 156144 465928 156196 465934
rect 156144 465870 156196 465876
rect 153384 465860 153436 465866
rect 153384 465802 153436 465808
rect 136088 465792 136140 465798
rect 136088 465734 136140 465740
rect 128728 465724 128780 465730
rect 128728 465666 128780 465672
rect 118608 465248 118660 465254
rect 91190 465216 91246 465225
rect 91190 465151 91246 465160
rect 96158 465216 96214 465225
rect 96158 465151 96214 465160
rect 98550 465216 98606 465225
rect 98550 465151 98606 465160
rect 101678 465216 101734 465225
rect 101678 465151 101734 465160
rect 103702 465216 103758 465225
rect 103702 465151 103758 465160
rect 111062 465216 111118 465225
rect 111062 465151 111118 465160
rect 113822 465216 113878 465225
rect 113822 465151 113878 465160
rect 116214 465216 116270 465225
rect 116214 465151 116216 465160
rect 116268 465151 116270 465160
rect 118606 465216 118608 465225
rect 128740 465225 128768 465666
rect 136100 465225 136128 465734
rect 153396 465225 153424 465802
rect 156156 465225 156184 465870
rect 168380 465656 168432 465662
rect 168380 465598 168432 465604
rect 168472 465656 168524 465662
rect 168472 465598 168524 465604
rect 118660 465216 118662 465225
rect 118606 465151 118662 465160
rect 128726 465216 128782 465225
rect 128726 465151 128782 465160
rect 136086 465216 136142 465225
rect 136086 465151 136142 465160
rect 141054 465216 141110 465225
rect 141054 465151 141110 465160
rect 143630 465216 143686 465225
rect 143630 465151 143686 465160
rect 153382 465216 153438 465225
rect 153382 465151 153438 465160
rect 156142 465216 156198 465225
rect 156142 465151 156198 465160
rect 116216 465122 116268 465128
rect 141068 465050 141096 465151
rect 143644 465118 143672 465151
rect 143632 465112 143684 465118
rect 143632 465054 143684 465060
rect 155868 465112 155920 465118
rect 155868 465054 155920 465060
rect 141056 465044 141108 465050
rect 141056 464986 141108 464992
rect 133512 464976 133564 464982
rect 133512 464918 133564 464924
rect 131120 464840 131172 464846
rect 131120 464782 131172 464788
rect 125968 464772 126020 464778
rect 125968 464714 126020 464720
rect 123576 464704 123628 464710
rect 123576 464646 123628 464652
rect 121000 464636 121052 464642
rect 121000 464578 121052 464584
rect 83464 464364 83516 464370
rect 83464 464306 83516 464312
rect 83476 463729 83504 464306
rect 121012 463729 121040 464578
rect 123588 463729 123616 464646
rect 125980 463729 126008 464714
rect 131132 464001 131160 464782
rect 131118 463992 131174 464001
rect 131118 463927 131174 463936
rect 133524 463729 133552 464918
rect 155880 464506 155908 465054
rect 168392 464574 168420 465598
rect 168484 465225 168512 465598
rect 169772 465225 169800 465938
rect 168470 465216 168526 465225
rect 168470 465151 168526 465160
rect 169758 465216 169814 465225
rect 169758 465151 169814 465160
rect 179432 464914 179460 465967
rect 186780 465928 186832 465934
rect 186780 465870 186832 465876
rect 186870 465896 186926 465905
rect 186688 465860 186740 465866
rect 186688 465802 186740 465808
rect 179420 464908 179472 464914
rect 179420 464850 179472 464856
rect 168380 464568 168432 464574
rect 168380 464510 168432 464516
rect 155868 464500 155920 464506
rect 155868 464442 155920 464448
rect 138480 464432 138532 464438
rect 138480 464374 138532 464380
rect 138492 463729 138520 464374
rect 146024 464296 146076 464302
rect 146024 464238 146076 464244
rect 146036 463729 146064 464238
rect 148508 464228 148560 464234
rect 148508 464170 148560 464176
rect 148520 463729 148548 464170
rect 151084 464160 151136 464166
rect 151084 464102 151136 464108
rect 151096 463729 151124 464102
rect 83462 463720 83518 463729
rect 83462 463655 83518 463664
rect 120998 463720 121054 463729
rect 120998 463655 121054 463664
rect 123574 463720 123630 463729
rect 123574 463655 123630 463664
rect 125966 463720 126022 463729
rect 125966 463655 126022 463664
rect 133510 463720 133566 463729
rect 133510 463655 133566 463664
rect 138478 463720 138534 463729
rect 138478 463655 138534 463664
rect 146022 463720 146078 463729
rect 146022 463655 146078 463664
rect 148506 463720 148562 463729
rect 148506 463655 148562 463664
rect 151082 463720 151138 463729
rect 151082 463655 151138 463664
rect 186700 463078 186728 465802
rect 186688 463072 186740 463078
rect 186688 463014 186740 463020
rect 186792 463010 186820 465870
rect 186870 465831 186926 465840
rect 186780 463004 186832 463010
rect 186780 462946 186832 462952
rect 186884 461553 186912 465831
rect 188342 465760 188398 465769
rect 187148 465724 187200 465730
rect 188342 465695 188398 465704
rect 187148 465666 187200 465672
rect 187056 464704 187108 464710
rect 187056 464646 187108 464652
rect 186964 464636 187016 464642
rect 186964 464578 187016 464584
rect 186870 461544 186926 461553
rect 186870 461479 186926 461488
rect 43444 448588 43496 448594
rect 43444 448530 43496 448536
rect 23480 181552 23532 181558
rect 23480 181494 23532 181500
rect 7562 179480 7618 179489
rect 7562 179415 7618 179424
rect 43456 179178 43484 448530
rect 48042 416936 48098 416945
rect 48042 416871 48098 416880
rect 47950 413808 48006 413817
rect 47950 413743 48006 413752
rect 46204 397520 46256 397526
rect 46204 397462 46256 397468
rect 46216 179246 46244 397462
rect 47582 388376 47638 388385
rect 47582 388311 47638 388320
rect 47596 207738 47624 388311
rect 47858 388104 47914 388113
rect 47858 388039 47914 388048
rect 47872 367810 47900 388039
rect 47964 378146 47992 413743
rect 47952 378140 48004 378146
rect 47952 378082 48004 378088
rect 47860 367804 47912 367810
rect 47860 367746 47912 367752
rect 48056 365702 48084 416871
rect 48134 415984 48190 415993
rect 48134 415919 48190 415928
rect 48044 365696 48096 365702
rect 48044 365638 48096 365644
rect 48148 359514 48176 415919
rect 49330 412856 49386 412865
rect 49330 412791 49386 412800
rect 49238 410000 49294 410009
rect 49238 409935 49294 409944
rect 48226 390008 48282 390017
rect 48226 389943 48282 389952
rect 48240 370530 48268 389943
rect 48228 370524 48280 370530
rect 48228 370466 48280 370472
rect 48136 359508 48188 359514
rect 48136 359450 48188 359456
rect 49252 313274 49280 409935
rect 49344 376038 49372 412791
rect 49422 411074 49478 411083
rect 49422 411009 49478 411018
rect 49332 376032 49384 376038
rect 49332 375974 49384 375980
rect 49436 347070 49464 411009
rect 49606 408218 49662 408227
rect 49606 408153 49662 408162
rect 49424 347064 49476 347070
rect 49424 347006 49476 347012
rect 49240 313268 49292 313274
rect 49240 313210 49292 313216
rect 49620 307766 49648 408153
rect 186688 380928 186740 380934
rect 186688 380870 186740 380876
rect 123482 379672 123538 379681
rect 123482 379607 123538 379616
rect 130934 379672 130990 379681
rect 130934 379607 130990 379616
rect 133510 379672 133566 379681
rect 133510 379607 133566 379616
rect 145930 379672 145986 379681
rect 145930 379607 145986 379616
rect 148506 379672 148562 379681
rect 148506 379607 148562 379616
rect 155958 379672 156014 379681
rect 155958 379607 156014 379616
rect 93950 379536 94006 379545
rect 93950 379471 94006 379480
rect 96434 379536 96490 379545
rect 96434 379471 96490 379480
rect 97630 379536 97686 379545
rect 97630 379471 97686 379480
rect 98734 379536 98790 379545
rect 98734 379471 98790 379480
rect 102230 379536 102286 379545
rect 102230 379471 102286 379480
rect 93964 378826 93992 379471
rect 96448 379098 96476 379471
rect 96436 379092 96488 379098
rect 96436 379034 96488 379040
rect 97644 378894 97672 379471
rect 98748 378962 98776 379471
rect 102244 379030 102272 379471
rect 123496 379234 123524 379607
rect 125966 379536 126022 379545
rect 125966 379471 126022 379480
rect 128542 379536 128598 379545
rect 128542 379471 128598 379480
rect 125980 379370 126008 379471
rect 125968 379364 126020 379370
rect 125968 379306 126020 379312
rect 128556 379302 128584 379471
rect 128544 379296 128596 379302
rect 128544 379238 128596 379244
rect 123484 379228 123536 379234
rect 123484 379170 123536 379176
rect 130948 379166 130976 379607
rect 133524 379438 133552 379607
rect 145944 379506 145972 379607
rect 145932 379500 145984 379506
rect 145932 379442 145984 379448
rect 133512 379432 133564 379438
rect 133512 379374 133564 379380
rect 130936 379160 130988 379166
rect 130936 379102 130988 379108
rect 102232 379024 102284 379030
rect 102232 378966 102284 378972
rect 98736 378956 98788 378962
rect 98736 378898 98788 378904
rect 97632 378888 97684 378894
rect 97632 378830 97684 378836
rect 93952 378820 94004 378826
rect 93952 378762 94004 378768
rect 148520 378758 148548 379607
rect 150990 379264 151046 379273
rect 150990 379199 151046 379208
rect 148508 378752 148560 378758
rect 148508 378694 148560 378700
rect 151004 378690 151032 379199
rect 150992 378684 151044 378690
rect 150992 378626 151044 378632
rect 155972 378622 156000 379607
rect 186700 379234 186728 380870
rect 186688 379228 186740 379234
rect 186688 379170 186740 379176
rect 155960 378616 156012 378622
rect 155960 378558 156012 378564
rect 50344 378140 50396 378146
rect 50344 378082 50396 378088
rect 95332 378140 95384 378146
rect 95332 378082 95384 378088
rect 50356 327078 50384 378082
rect 95344 378049 95372 378082
rect 99840 378072 99892 378078
rect 67546 378040 67602 378049
rect 67546 377975 67602 377984
rect 73158 378040 73214 378049
rect 73158 377975 73214 377984
rect 74354 378040 74410 378049
rect 74354 377975 74410 377984
rect 78494 378040 78550 378049
rect 78494 377975 78550 377984
rect 81162 378040 81218 378049
rect 81162 377975 81218 377984
rect 92294 378040 92350 378049
rect 92294 377975 92350 377984
rect 92846 378040 92902 378049
rect 92846 377975 92902 377984
rect 95330 378040 95386 378049
rect 95330 377975 95386 377984
rect 96526 378040 96582 378049
rect 96526 377975 96582 377984
rect 99838 378040 99840 378049
rect 99892 378040 99894 378049
rect 99838 377975 99894 377984
rect 101310 378040 101366 378049
rect 101310 377975 101312 377984
rect 66166 377088 66222 377097
rect 66166 377023 66222 377032
rect 50436 365696 50488 365702
rect 50436 365638 50488 365644
rect 50448 335306 50476 365638
rect 50436 335300 50488 335306
rect 50436 335242 50488 335248
rect 50344 327072 50396 327078
rect 50344 327014 50396 327020
rect 49608 307760 49660 307766
rect 49608 307702 49660 307708
rect 66180 296682 66208 377023
rect 67560 302190 67588 377975
rect 73172 377874 73200 377975
rect 73160 377868 73212 377874
rect 73160 377810 73212 377816
rect 68926 377088 68982 377097
rect 68926 377023 68982 377032
rect 70306 377088 70362 377097
rect 70306 377023 70362 377032
rect 71686 377088 71742 377097
rect 71686 377023 71742 377032
rect 73066 377088 73122 377097
rect 73066 377023 73122 377032
rect 67548 302184 67600 302190
rect 67548 302126 67600 302132
rect 68940 300830 68968 377023
rect 70320 306338 70348 377023
rect 71700 311846 71728 377023
rect 73080 317422 73108 377023
rect 73068 317416 73120 317422
rect 73068 317358 73120 317364
rect 71688 311840 71740 311846
rect 71688 311782 71740 311788
rect 70308 306332 70360 306338
rect 70308 306274 70360 306280
rect 74368 303618 74396 377975
rect 75184 377868 75236 377874
rect 75184 377810 75236 377816
rect 74356 303612 74408 303618
rect 74356 303554 74408 303560
rect 68928 300824 68980 300830
rect 68928 300766 68980 300772
rect 75196 299470 75224 377810
rect 75826 377088 75882 377097
rect 75826 377023 75882 377032
rect 77206 377088 77262 377097
rect 77206 377023 77262 377032
rect 78310 377088 78366 377097
rect 78310 377023 78312 377032
rect 75840 309126 75868 377023
rect 77220 314634 77248 377023
rect 78364 377023 78366 377032
rect 78312 376994 78364 377000
rect 78508 320142 78536 377975
rect 79966 377088 80022 377097
rect 79324 377052 79376 377058
rect 79966 377023 80022 377032
rect 79324 376994 79376 377000
rect 78496 320136 78548 320142
rect 78496 320078 78548 320084
rect 77208 314628 77260 314634
rect 77208 314570 77260 314576
rect 75828 309120 75880 309126
rect 75828 309062 75880 309068
rect 75184 299464 75236 299470
rect 75184 299406 75236 299412
rect 79336 299402 79364 376994
rect 79980 324290 80008 377023
rect 81176 332586 81204 377975
rect 81254 377088 81310 377097
rect 81254 377023 81310 377032
rect 82726 377088 82782 377097
rect 82726 377023 82782 377032
rect 84106 377088 84162 377097
rect 84106 377023 84162 377032
rect 85486 377088 85542 377097
rect 85486 377023 85542 377032
rect 86866 377088 86922 377097
rect 86866 377023 86922 377032
rect 88154 377088 88210 377097
rect 88154 377023 88210 377032
rect 89534 377088 89590 377097
rect 89534 377023 89590 377032
rect 91006 377088 91062 377097
rect 91006 377023 91062 377032
rect 91742 377088 91798 377097
rect 91742 377023 91744 377032
rect 81164 332580 81216 332586
rect 81164 332522 81216 332528
rect 81268 328438 81296 377023
rect 81346 376952 81402 376961
rect 81346 376887 81402 376896
rect 81256 328432 81308 328438
rect 81256 328374 81308 328380
rect 79968 324284 80020 324290
rect 79968 324226 80020 324232
rect 81360 304978 81388 376887
rect 82740 338094 82768 377023
rect 84014 376952 84070 376961
rect 84014 376887 84070 376896
rect 84028 342242 84056 376887
rect 84016 342236 84068 342242
rect 84016 342178 84068 342184
rect 82728 338088 82780 338094
rect 82728 338030 82780 338036
rect 84120 310486 84148 377023
rect 85500 346390 85528 377023
rect 86774 376952 86830 376961
rect 86774 376887 86830 376896
rect 86788 350538 86816 376887
rect 86776 350532 86828 350538
rect 86776 350474 86828 350480
rect 85488 346384 85540 346390
rect 85488 346326 85540 346332
rect 86880 315994 86908 377023
rect 88168 358766 88196 377023
rect 88246 376952 88302 376961
rect 88246 376887 88302 376896
rect 88156 358760 88208 358766
rect 88156 358702 88208 358708
rect 88260 354686 88288 376887
rect 89548 364342 89576 377023
rect 89626 376952 89682 376961
rect 89626 376887 89682 376896
rect 89536 364336 89588 364342
rect 89536 364278 89588 364284
rect 88248 354680 88300 354686
rect 88248 354622 88300 354628
rect 89640 320074 89668 376887
rect 91020 368490 91048 377023
rect 91796 377023 91798 377032
rect 91744 376994 91796 377000
rect 92308 372570 92336 377975
rect 92860 376718 92888 377975
rect 93766 377088 93822 377097
rect 93124 377052 93176 377058
rect 93766 377023 93822 377032
rect 93124 376994 93176 377000
rect 92848 376712 92900 376718
rect 92848 376654 92900 376660
rect 92296 372564 92348 372570
rect 92296 372506 92348 372512
rect 91008 368484 91060 368490
rect 91008 368426 91060 368432
rect 93136 325650 93164 376994
rect 93780 329798 93808 377023
rect 96540 333946 96568 377975
rect 101364 377975 101366 377984
rect 103334 378040 103390 378049
rect 103334 377975 103390 377984
rect 104806 378040 104862 378049
rect 104806 377975 104862 377984
rect 105910 378040 105966 378049
rect 105910 377975 105966 377984
rect 107566 378040 107622 378049
rect 107566 377975 107622 377984
rect 110234 378040 110290 378049
rect 110234 377975 110290 377984
rect 114466 378040 114522 378049
rect 114466 377975 114522 377984
rect 120998 378040 121054 378049
rect 120998 377975 121054 377984
rect 136086 378040 136142 378049
rect 136086 377975 136142 377984
rect 139030 378040 139086 378049
rect 139030 377975 139086 377984
rect 141606 378040 141662 378049
rect 141606 377975 141662 377984
rect 143446 378040 143502 378049
rect 143446 377975 143502 377984
rect 153382 378040 153438 378049
rect 153382 377975 153438 377984
rect 101312 377946 101364 377952
rect 103348 377942 103376 377975
rect 103336 377936 103388 377942
rect 103336 377878 103388 377884
rect 104438 377904 104494 377913
rect 104438 377839 104440 377848
rect 104492 377839 104494 377848
rect 104440 377810 104492 377816
rect 99286 377088 99342 377097
rect 99286 377023 99342 377032
rect 102046 377088 102102 377097
rect 102046 377023 102102 377032
rect 99300 338026 99328 377023
rect 102060 342174 102088 377023
rect 104820 347750 104848 377975
rect 105924 377738 105952 377975
rect 107580 377806 107608 377975
rect 107568 377800 107620 377806
rect 107568 377742 107620 377748
rect 105912 377732 105964 377738
rect 105912 377674 105964 377680
rect 110248 377670 110276 377975
rect 110236 377664 110288 377670
rect 110236 377606 110288 377612
rect 106186 377088 106242 377097
rect 106186 377023 106242 377032
rect 108946 377088 109002 377097
rect 108946 377023 109002 377032
rect 111706 377088 111762 377097
rect 111706 377023 111762 377032
rect 106200 351898 106228 377023
rect 108960 356046 108988 377023
rect 111720 360194 111748 377023
rect 114480 364274 114508 377975
rect 121012 377466 121040 377975
rect 136100 377602 136128 377975
rect 136088 377596 136140 377602
rect 136088 377538 136140 377544
rect 139044 377534 139072 377975
rect 139032 377528 139084 377534
rect 139032 377470 139084 377476
rect 121000 377460 121052 377466
rect 121000 377402 121052 377408
rect 141620 377398 141648 377975
rect 141608 377392 141660 377398
rect 141608 377334 141660 377340
rect 143460 377330 143488 377975
rect 143448 377324 143500 377330
rect 143448 377266 143500 377272
rect 153396 377262 153424 377975
rect 180706 377360 180762 377369
rect 180706 377295 180762 377304
rect 153384 377256 153436 377262
rect 153384 377198 153436 377204
rect 117226 377088 117282 377097
rect 117226 377023 117282 377032
rect 118606 377088 118662 377097
rect 118606 377023 118662 377032
rect 173714 377088 173770 377097
rect 173714 377023 173770 377032
rect 117240 368422 117268 377023
rect 118620 373998 118648 377023
rect 118608 373992 118660 373998
rect 118608 373934 118660 373940
rect 148324 370524 148376 370530
rect 148324 370466 148376 370472
rect 117228 368416 117280 368422
rect 117228 368358 117280 368364
rect 122104 367804 122156 367810
rect 122104 367746 122156 367752
rect 114468 364268 114520 364274
rect 114468 364210 114520 364216
rect 111708 360188 111760 360194
rect 111708 360130 111760 360136
rect 108948 356040 109000 356046
rect 108948 355982 109000 355988
rect 106188 351892 106240 351898
rect 106188 351834 106240 351840
rect 104808 347744 104860 347750
rect 104808 347686 104860 347692
rect 102048 342168 102100 342174
rect 102048 342110 102100 342116
rect 99288 338020 99340 338026
rect 99288 337962 99340 337968
rect 96528 333940 96580 333946
rect 96528 333882 96580 333888
rect 93768 329792 93820 329798
rect 93768 329734 93820 329740
rect 93124 325644 93176 325650
rect 93124 325586 93176 325592
rect 89628 320068 89680 320074
rect 89628 320010 89680 320016
rect 86868 315988 86920 315994
rect 86868 315930 86920 315936
rect 84108 310480 84160 310486
rect 84108 310422 84160 310428
rect 81348 304972 81400 304978
rect 81348 304914 81400 304920
rect 79324 299396 79376 299402
rect 79324 299338 79376 299344
rect 66168 296676 66220 296682
rect 66168 296618 66220 296624
rect 122116 293962 122144 367746
rect 148336 296614 148364 370466
rect 167644 359508 167696 359514
rect 167644 359450 167696 359456
rect 167656 331226 167684 359450
rect 173728 336734 173756 377023
rect 173806 376952 173862 376961
rect 173806 376887 173862 376896
rect 173716 336728 173768 336734
rect 173716 336670 173768 336676
rect 173820 332518 173848 376887
rect 173808 332512 173860 332518
rect 173808 332454 173860 332460
rect 167644 331220 167696 331226
rect 167644 331162 167696 331168
rect 148324 296608 148376 296614
rect 148324 296550 148376 296556
rect 122104 293956 122156 293962
rect 122104 293898 122156 293904
rect 157248 292664 157300 292670
rect 157248 292606 157300 292612
rect 154488 289876 154540 289882
rect 154488 289818 154540 289824
rect 151728 287088 151780 287094
rect 151728 287030 151780 287036
rect 144828 286476 144880 286482
rect 144828 286418 144880 286424
rect 141884 286408 141936 286414
rect 49606 286376 49662 286385
rect 141884 286350 141936 286356
rect 49606 286311 49662 286320
rect 139308 286340 139360 286346
rect 48134 236872 48190 236881
rect 48134 236807 48190 236816
rect 47950 235920 48006 235929
rect 47950 235855 48006 235864
rect 47858 233744 47914 233753
rect 47858 233679 47914 233688
rect 47766 231024 47822 231033
rect 47766 230959 47822 230968
rect 47674 229936 47730 229945
rect 47674 229871 47730 229880
rect 47584 207732 47636 207738
rect 47584 207674 47636 207680
rect 47688 199073 47716 229871
rect 47674 199064 47730 199073
rect 47674 198999 47730 199008
rect 47780 197198 47808 230959
rect 47872 199753 47900 233679
rect 47964 199889 47992 235855
rect 48042 232792 48098 232801
rect 48042 232727 48098 232736
rect 47950 199880 48006 199889
rect 47950 199815 48006 199824
rect 47858 199744 47914 199753
rect 47858 199679 47914 199688
rect 47768 197192 47820 197198
rect 47768 197134 47820 197140
rect 48056 197130 48084 232727
rect 48148 199617 48176 236807
rect 49514 228218 49570 228227
rect 49514 228153 49570 228162
rect 49330 209944 49386 209953
rect 49330 209879 49386 209888
rect 48228 207732 48280 207738
rect 48228 207674 48280 207680
rect 48134 199608 48190 199617
rect 48134 199543 48190 199552
rect 48044 197124 48096 197130
rect 48044 197066 48096 197072
rect 48240 182714 48268 207674
rect 47584 182708 47636 182714
rect 47584 182650 47636 182656
rect 48228 182708 48280 182714
rect 48228 182650 48280 182656
rect 46204 179240 46256 179246
rect 46204 179182 46256 179188
rect 43444 179172 43496 179178
rect 43444 179114 43496 179120
rect 6184 176656 6236 176662
rect 6184 176598 6236 176604
rect 3424 150408 3476 150414
rect 3424 150350 3476 150356
rect 3436 149841 3464 150350
rect 3422 149832 3478 149841
rect 3422 149767 3478 149776
rect 3332 141432 3384 141438
rect 3332 141374 3384 141380
rect 3344 136785 3372 141374
rect 3330 136776 3386 136785
rect 3330 136711 3386 136720
rect 3148 85536 3200 85542
rect 3148 85478 3200 85484
rect 3160 84697 3188 85478
rect 3146 84688 3202 84697
rect 3146 84623 3202 84632
rect 3424 45552 3476 45558
rect 3422 45520 3424 45529
rect 3476 45520 3478 45529
rect 3422 45455 3478 45464
rect 3424 6860 3476 6866
rect 3424 6802 3476 6808
rect 3436 6497 3464 6802
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 47596 3466 47624 182650
rect 48240 182238 48268 182650
rect 48228 182232 48280 182238
rect 48228 182174 48280 182180
rect 49344 182170 49372 209879
rect 49422 208090 49478 208099
rect 49422 208025 49478 208034
rect 49436 182850 49464 208025
rect 49528 194546 49556 228153
rect 49620 208371 49648 286311
rect 139308 286282 139360 286288
rect 136548 286272 136600 286278
rect 136546 286240 136548 286249
rect 139320 286249 139348 286282
rect 136600 286240 136602 286249
rect 126888 286204 126940 286210
rect 136546 286175 136602 286184
rect 139306 286240 139362 286249
rect 139306 286175 139362 286184
rect 126888 286146 126940 286152
rect 124128 286136 124180 286142
rect 124128 286078 124180 286084
rect 108948 286068 109000 286074
rect 108948 286010 109000 286016
rect 106188 286000 106240 286006
rect 106186 285968 106188 285977
rect 108960 285977 108988 286010
rect 106240 285968 106242 285977
rect 104808 285932 104860 285938
rect 106186 285903 106242 285912
rect 108946 285968 109002 285977
rect 108946 285903 109002 285912
rect 104808 285874 104860 285880
rect 83740 285728 83792 285734
rect 83738 285696 83740 285705
rect 104820 285705 104848 285874
rect 118608 285864 118660 285870
rect 118608 285806 118660 285812
rect 114468 285796 114520 285802
rect 114468 285738 114520 285744
rect 114480 285705 114508 285738
rect 118620 285705 118648 285806
rect 124140 285705 124168 286078
rect 126900 285705 126928 286146
rect 141896 285705 141924 286350
rect 144840 286249 144868 286418
rect 144826 286240 144882 286249
rect 144826 286175 144882 286184
rect 151740 285705 151768 287030
rect 154500 285705 154528 289818
rect 157260 285705 157288 292606
rect 170680 286612 170732 286618
rect 170680 286554 170732 286560
rect 169668 286544 169720 286550
rect 169668 286486 169720 286492
rect 169680 285705 169708 286486
rect 170692 286249 170720 286554
rect 180720 286385 180748 377295
rect 186976 376961 187004 464578
rect 187068 383654 187096 464646
rect 187160 391950 187188 465666
rect 187698 465216 187754 465225
rect 187698 465151 187754 465160
rect 187148 391944 187200 391950
rect 187148 391886 187200 391892
rect 187056 383648 187108 383654
rect 187056 383590 187108 383596
rect 187712 377369 187740 465151
rect 188160 385076 188212 385082
rect 188160 385018 188212 385024
rect 188172 379370 188200 385018
rect 188160 379364 188212 379370
rect 188160 379306 188212 379312
rect 187698 377360 187754 377369
rect 187698 377295 187754 377304
rect 186962 376952 187018 376961
rect 186962 376887 187018 376896
rect 188356 306270 188384 465695
rect 188436 465588 188488 465594
rect 188436 465530 188488 465536
rect 188448 361554 188476 465530
rect 189724 465520 189776 465526
rect 189724 465462 189776 465468
rect 188712 464976 188764 464982
rect 188712 464918 188764 464924
rect 188620 464840 188672 464846
rect 188620 464782 188672 464788
rect 188528 464772 188580 464778
rect 188528 464714 188580 464720
rect 188540 387802 188568 464714
rect 188632 396030 188660 464782
rect 188724 400178 188752 464918
rect 189078 459232 189134 459241
rect 189078 459167 189134 459176
rect 189092 458250 189120 459167
rect 189080 458244 189132 458250
rect 189080 458186 189132 458192
rect 188804 433356 188856 433362
rect 188804 433298 188856 433304
rect 188712 400172 188764 400178
rect 188712 400114 188764 400120
rect 188620 396024 188672 396030
rect 188620 395966 188672 395972
rect 188528 387796 188580 387802
rect 188528 387738 188580 387744
rect 188816 377262 188844 433298
rect 189078 399392 189134 399401
rect 189078 399327 189134 399336
rect 189092 398886 189120 399327
rect 189080 398880 189132 398886
rect 189080 398822 189132 398828
rect 189078 397760 189134 397769
rect 189078 397695 189134 397704
rect 189092 397526 189120 397695
rect 189080 397520 189132 397526
rect 189080 397462 189132 397468
rect 189262 396400 189318 396409
rect 189262 396335 189318 396344
rect 189276 396098 189304 396335
rect 189264 396092 189316 396098
rect 189264 396034 189316 396040
rect 189078 394904 189134 394913
rect 189078 394839 189134 394848
rect 189092 394738 189120 394839
rect 189080 394732 189132 394738
rect 189080 394674 189132 394680
rect 189262 393680 189318 393689
rect 189262 393615 189318 393624
rect 189276 393378 189304 393615
rect 189264 393372 189316 393378
rect 189264 393314 189316 393320
rect 188804 377256 188856 377262
rect 188804 377198 188856 377204
rect 188436 361548 188488 361554
rect 188436 361490 188488 361496
rect 189736 343602 189764 465462
rect 189908 464160 189960 464166
rect 189908 464102 189960 464108
rect 189816 437504 189868 437510
rect 189816 437446 189868 437452
rect 189828 377670 189856 437446
rect 189920 431934 189948 464102
rect 189908 431928 189960 431934
rect 189908 431870 189960 431876
rect 189908 389224 189960 389230
rect 189908 389166 189960 389172
rect 189920 379098 189948 389166
rect 189908 379092 189960 379098
rect 189908 379034 189960 379040
rect 189816 377664 189868 377670
rect 189816 377606 189868 377612
rect 189724 343596 189776 343602
rect 189724 343538 189776 343544
rect 188344 306264 188396 306270
rect 188344 306206 188396 306212
rect 186780 286476 186832 286482
rect 186780 286418 186832 286424
rect 180706 286376 180762 286385
rect 180706 286311 180762 286320
rect 170678 286240 170734 286249
rect 170678 286175 170734 286184
rect 83792 285696 83794 285705
rect 83738 285631 83794 285640
rect 86866 285696 86922 285705
rect 86866 285631 86922 285640
rect 89626 285696 89682 285705
rect 89626 285631 89682 285640
rect 92386 285696 92442 285705
rect 92386 285631 92388 285640
rect 86880 285462 86908 285631
rect 86868 285456 86920 285462
rect 86868 285398 86920 285404
rect 89640 285326 89668 285631
rect 92440 285631 92442 285640
rect 93674 285696 93730 285705
rect 93674 285631 93730 285640
rect 96526 285696 96582 285705
rect 96526 285631 96582 285640
rect 104806 285696 104862 285705
rect 104806 285631 104862 285640
rect 114466 285696 114522 285705
rect 114466 285631 114522 285640
rect 118606 285696 118662 285705
rect 118606 285631 118662 285640
rect 124126 285696 124182 285705
rect 124126 285631 124182 285640
rect 126886 285696 126942 285705
rect 126886 285631 126942 285640
rect 133786 285696 133842 285705
rect 133786 285631 133842 285640
rect 141882 285696 141938 285705
rect 141882 285631 141938 285640
rect 151726 285696 151782 285705
rect 151726 285631 151782 285640
rect 154486 285696 154542 285705
rect 154486 285631 154542 285640
rect 157246 285696 157302 285705
rect 157246 285631 157302 285640
rect 169666 285696 169722 285705
rect 169666 285631 169722 285640
rect 92388 285602 92440 285608
rect 93688 285598 93716 285631
rect 93676 285592 93728 285598
rect 93676 285534 93728 285540
rect 96540 285530 96568 285631
rect 96528 285524 96580 285530
rect 96528 285466 96580 285472
rect 133800 285394 133828 285631
rect 133788 285388 133840 285394
rect 133788 285330 133840 285336
rect 89628 285320 89680 285326
rect 89628 285262 89680 285268
rect 131120 285252 131172 285258
rect 131120 285194 131172 285200
rect 128728 285184 128780 285190
rect 128726 285152 128728 285161
rect 131132 285161 131160 285194
rect 128780 285152 128782 285161
rect 116216 285116 116268 285122
rect 128726 285087 128782 285096
rect 131118 285152 131174 285161
rect 131118 285087 131174 285096
rect 116216 285058 116268 285064
rect 111064 285048 111116 285054
rect 111062 285016 111064 285025
rect 116228 285025 116256 285058
rect 111116 285016 111118 285025
rect 98552 284980 98604 284986
rect 111062 284951 111118 284960
rect 116214 285016 116270 285025
rect 116214 284951 116270 284960
rect 98552 284922 98604 284928
rect 98564 284889 98592 284922
rect 148600 284912 148652 284918
rect 98550 284880 98606 284889
rect 148598 284880 148600 284889
rect 148652 284880 148654 284889
rect 98550 284815 98606 284824
rect 101312 284844 101364 284850
rect 148598 284815 148654 284824
rect 101312 284786 101364 284792
rect 101324 284753 101352 284786
rect 146024 284776 146076 284782
rect 101310 284744 101366 284753
rect 101310 284679 101366 284688
rect 146022 284744 146024 284753
rect 146076 284744 146078 284753
rect 146022 284679 146078 284688
rect 180720 284073 180748 286311
rect 186688 284776 186740 284782
rect 186688 284718 186740 284724
rect 180706 284064 180762 284073
rect 180706 283999 180762 284008
rect 186700 282878 186728 284718
rect 186688 282872 186740 282878
rect 186688 282814 186740 282820
rect 186792 280158 186820 286418
rect 187332 286408 187384 286414
rect 187332 286350 187384 286356
rect 187240 286340 187292 286346
rect 187240 286282 187292 286288
rect 187148 286272 187200 286278
rect 187148 286214 187200 286220
rect 187056 286204 187108 286210
rect 187056 286146 187108 286152
rect 186964 286136 187016 286142
rect 186964 286078 187016 286084
rect 186780 280152 186832 280158
rect 186780 280094 186832 280100
rect 186976 259418 187004 286078
rect 187068 262206 187096 286146
rect 187160 271862 187188 286214
rect 187252 274650 187280 286282
rect 187344 277370 187372 286350
rect 189724 285456 189776 285462
rect 189724 285398 189776 285404
rect 187608 280220 187660 280226
rect 187608 280162 187660 280168
rect 187332 277364 187384 277370
rect 187332 277306 187384 277312
rect 187240 274644 187292 274650
rect 187240 274586 187292 274592
rect 187148 271856 187200 271862
rect 187148 271798 187200 271804
rect 187056 262200 187108 262206
rect 187056 262142 187108 262148
rect 187148 260908 187200 260914
rect 187148 260850 187200 260856
rect 186964 259412 187016 259418
rect 186964 259354 187016 259360
rect 186964 241528 187016 241534
rect 186964 241470 187016 241476
rect 49606 208362 49662 208371
rect 49606 208297 49662 208306
rect 49620 207738 49648 208297
rect 49608 207732 49660 207738
rect 49608 207674 49660 207680
rect 136548 199572 136600 199578
rect 136548 199514 136600 199520
rect 106004 199504 106056 199510
rect 71870 199472 71926 199481
rect 71870 199407 71926 199416
rect 77758 199472 77814 199481
rect 77758 199407 77814 199416
rect 81346 199472 81402 199481
rect 81346 199407 81402 199416
rect 82542 199472 82598 199481
rect 82542 199407 82598 199416
rect 83462 199472 83518 199481
rect 83462 199407 83518 199416
rect 86222 199472 86278 199481
rect 86222 199407 86278 199416
rect 103702 199472 103758 199481
rect 106004 199446 106056 199452
rect 103702 199407 103704 199416
rect 71884 198966 71912 199407
rect 77772 199034 77800 199407
rect 81360 199102 81388 199407
rect 82556 199170 82584 199407
rect 83476 199238 83504 199407
rect 86236 199306 86264 199407
rect 103756 199407 103758 199416
rect 103704 199378 103756 199384
rect 86224 199300 86276 199306
rect 86224 199242 86276 199248
rect 83464 199232 83516 199238
rect 83464 199174 83516 199180
rect 82544 199164 82596 199170
rect 82544 199106 82596 199112
rect 81348 199096 81400 199102
rect 81348 199038 81400 199044
rect 77760 199028 77812 199034
rect 77760 198970 77812 198976
rect 71872 198960 71924 198966
rect 71872 198902 71924 198908
rect 91192 198892 91244 198898
rect 91192 198834 91244 198840
rect 88616 198824 88668 198830
rect 88616 198766 88668 198772
rect 78864 198756 78916 198762
rect 78864 198698 78916 198704
rect 78876 198665 78904 198698
rect 84568 198688 84620 198694
rect 70582 198656 70638 198665
rect 70582 198591 70638 198600
rect 76654 198656 76710 198665
rect 76654 198591 76710 198600
rect 78862 198656 78918 198665
rect 78862 198591 78918 198600
rect 80150 198656 80206 198665
rect 80150 198591 80206 198600
rect 84566 198656 84568 198665
rect 88628 198665 88656 198766
rect 91204 198665 91232 198834
rect 84620 198656 84622 198665
rect 84566 198591 84622 198600
rect 88246 198656 88302 198665
rect 88246 198591 88248 198600
rect 67546 198248 67602 198257
rect 67546 198183 67602 198192
rect 66166 197432 66222 197441
rect 66166 197367 66222 197376
rect 49516 194540 49568 194546
rect 49516 194482 49568 194488
rect 66180 183530 66208 197367
rect 67560 189038 67588 198183
rect 70596 198014 70624 198591
rect 74354 198248 74410 198257
rect 76668 198218 76696 198591
rect 80164 198422 80192 198591
rect 88300 198591 88302 198600
rect 88614 198656 88670 198665
rect 88614 198591 88670 198600
rect 91190 198656 91246 198665
rect 91190 198591 91246 198600
rect 93582 198656 93638 198665
rect 93582 198591 93638 198600
rect 93950 198656 94006 198665
rect 93950 198591 94006 198600
rect 95974 198656 96030 198665
rect 95974 198591 96030 198600
rect 98366 198656 98422 198665
rect 98366 198591 98422 198600
rect 99838 198656 99894 198665
rect 99838 198591 99894 198600
rect 100942 198656 100998 198665
rect 100942 198591 100998 198600
rect 102230 198656 102286 198665
rect 102230 198591 102286 198600
rect 88248 198562 88300 198568
rect 93596 198558 93624 198591
rect 93584 198552 93636 198558
rect 85854 198520 85910 198529
rect 85854 198455 85910 198464
rect 87418 198520 87474 198529
rect 87418 198455 87474 198464
rect 90914 198520 90970 198529
rect 93584 198494 93636 198500
rect 93964 198490 93992 198591
rect 90914 198455 90970 198464
rect 93952 198484 94004 198490
rect 80152 198416 80204 198422
rect 80152 198358 80204 198364
rect 74354 198183 74410 198192
rect 76656 198212 76708 198218
rect 70584 198008 70636 198014
rect 70584 197950 70636 197956
rect 68926 197432 68982 197441
rect 68926 197367 68982 197376
rect 69846 197432 69902 197441
rect 69846 197367 69902 197376
rect 67548 189032 67600 189038
rect 67548 188974 67600 188980
rect 68940 187678 68968 197367
rect 69860 193186 69888 197367
rect 69848 193180 69900 193186
rect 69848 193122 69900 193128
rect 74368 190466 74396 198183
rect 76656 198154 76708 198160
rect 75734 198112 75790 198121
rect 75734 198047 75790 198056
rect 74446 197432 74502 197441
rect 74446 197367 74502 197376
rect 74356 190460 74408 190466
rect 74356 190402 74408 190408
rect 68928 187672 68980 187678
rect 68928 187614 68980 187620
rect 74460 184890 74488 197367
rect 75748 195974 75776 198047
rect 83738 197976 83794 197985
rect 83738 197911 83794 197920
rect 78586 197432 78642 197441
rect 78586 197367 78642 197376
rect 81070 197432 81126 197441
rect 81070 197367 81126 197376
rect 75736 195968 75788 195974
rect 75736 195910 75788 195916
rect 78600 186318 78628 197367
rect 81084 191826 81112 197367
rect 83752 195906 83780 197911
rect 85868 196926 85896 198455
rect 85856 196920 85908 196926
rect 85856 196862 85908 196868
rect 87432 196858 87460 198455
rect 89534 198384 89590 198393
rect 89534 198319 89590 198328
rect 87420 196852 87472 196858
rect 87420 196794 87472 196800
rect 89548 196518 89576 198319
rect 90928 196790 90956 198455
rect 93952 198426 94004 198432
rect 92846 198384 92902 198393
rect 95988 198354 96016 198591
rect 92846 198319 92902 198328
rect 95976 198348 96028 198354
rect 92294 198248 92350 198257
rect 92294 198183 92350 198192
rect 90916 196784 90968 196790
rect 90916 196726 90968 196732
rect 89536 196512 89588 196518
rect 89536 196454 89588 196460
rect 92308 196450 92336 198183
rect 92860 196722 92888 198319
rect 95976 198290 96028 198296
rect 98380 198286 98408 198591
rect 98368 198280 98420 198286
rect 98368 198222 98420 198228
rect 99852 197946 99880 198591
rect 100956 198150 100984 198591
rect 100944 198144 100996 198150
rect 100944 198086 100996 198092
rect 99840 197940 99892 197946
rect 99840 197882 99892 197888
rect 92848 196716 92900 196722
rect 92848 196658 92900 196664
rect 102244 196654 102272 198591
rect 106016 198422 106044 199446
rect 128358 199336 128414 199345
rect 128358 199271 128414 199280
rect 106094 198656 106150 198665
rect 106094 198591 106150 198600
rect 107014 198656 107070 198665
rect 107014 198591 107070 198600
rect 108486 198656 108542 198665
rect 108486 198591 108542 198600
rect 113638 198656 113694 198665
rect 113638 198591 113694 198600
rect 120998 198656 121054 198665
rect 120998 198591 121054 198600
rect 123574 198656 123630 198665
rect 123574 198591 123630 198600
rect 106108 198422 106136 198591
rect 106004 198416 106056 198422
rect 106004 198358 106056 198364
rect 106096 198416 106148 198422
rect 106096 198358 106148 198364
rect 105910 197976 105966 197985
rect 105910 197911 105966 197920
rect 105924 197062 105952 197911
rect 105912 197056 105964 197062
rect 105912 196998 105964 197004
rect 107028 196994 107056 198591
rect 107016 196988 107068 196994
rect 107016 196930 107068 196936
rect 102232 196648 102284 196654
rect 102232 196590 102284 196596
rect 108500 196586 108528 198591
rect 111062 197976 111118 197985
rect 111062 197911 111118 197920
rect 108488 196580 108540 196586
rect 108488 196522 108540 196528
rect 92296 196444 92348 196450
rect 92296 196386 92348 196392
rect 83740 195900 83792 195906
rect 83740 195842 83792 195848
rect 111076 195838 111104 197911
rect 111064 195832 111116 195838
rect 111064 195774 111116 195780
rect 113652 195770 113680 198591
rect 116214 197840 116270 197849
rect 116214 197775 116270 197784
rect 118422 197840 118478 197849
rect 118422 197775 118478 197784
rect 113640 195764 113692 195770
rect 113640 195706 113692 195712
rect 116228 195634 116256 197775
rect 116216 195628 116268 195634
rect 116216 195570 116268 195576
rect 118436 195498 118464 197775
rect 118424 195492 118476 195498
rect 118424 195434 118476 195440
rect 121012 195430 121040 198591
rect 123588 198082 123616 198591
rect 123576 198076 123628 198082
rect 123576 198018 123628 198024
rect 128372 197946 128400 199271
rect 128542 198656 128598 198665
rect 128542 198591 128598 198600
rect 130934 198656 130990 198665
rect 130934 198591 130990 198600
rect 136086 198656 136142 198665
rect 136086 198591 136142 198600
rect 128556 197946 128584 198591
rect 128360 197940 128412 197946
rect 128360 197882 128412 197888
rect 128544 197940 128596 197946
rect 128544 197882 128596 197888
rect 130948 197878 130976 198591
rect 130936 197872 130988 197878
rect 130936 197814 130988 197820
rect 136100 197810 136128 198591
rect 136560 198218 136588 199514
rect 150990 199472 151046 199481
rect 150990 199407 151046 199416
rect 151004 199374 151032 199407
rect 150992 199368 151044 199374
rect 150992 199310 151044 199316
rect 138754 198656 138810 198665
rect 138754 198591 138810 198600
rect 143446 198656 143502 198665
rect 143446 198591 143502 198600
rect 146022 198656 146078 198665
rect 146022 198591 146078 198600
rect 148598 198656 148654 198665
rect 148598 198591 148654 198600
rect 153382 198656 153438 198665
rect 153382 198591 153438 198600
rect 173438 198656 173494 198665
rect 173438 198591 173494 198600
rect 136548 198212 136600 198218
rect 136548 198154 136600 198160
rect 136088 197804 136140 197810
rect 136088 197746 136140 197752
rect 126150 197704 126206 197713
rect 126150 197639 126206 197648
rect 133510 197704 133566 197713
rect 133510 197639 133566 197648
rect 121000 195424 121052 195430
rect 121000 195366 121052 195372
rect 126164 195362 126192 197639
rect 126152 195356 126204 195362
rect 126152 195298 126204 195304
rect 133524 195294 133552 197639
rect 138768 196897 138796 198591
rect 138754 196888 138810 196897
rect 138754 196823 138810 196832
rect 143460 196761 143488 198591
rect 143446 196752 143502 196761
rect 143446 196687 143502 196696
rect 133512 195288 133564 195294
rect 133512 195230 133564 195236
rect 146036 195226 146064 198591
rect 148612 198218 148640 198591
rect 148600 198212 148652 198218
rect 148600 198154 148652 198160
rect 153396 195702 153424 198591
rect 155958 197840 156014 197849
rect 155958 197775 156014 197784
rect 173254 197840 173310 197849
rect 173254 197775 173310 197784
rect 153384 195696 153436 195702
rect 153384 195638 153436 195644
rect 155972 195566 156000 197775
rect 173268 197266 173296 197775
rect 173452 197334 173480 198591
rect 173440 197328 173492 197334
rect 173440 197270 173492 197276
rect 173256 197260 173308 197266
rect 173256 197202 173308 197208
rect 186976 196586 187004 241470
rect 187056 227792 187108 227798
rect 187056 227734 187108 227740
rect 187068 199238 187096 227734
rect 187056 199232 187108 199238
rect 187056 199174 187108 199180
rect 187160 198529 187188 260850
rect 187332 259480 187384 259486
rect 187332 259422 187384 259428
rect 187240 222216 187292 222222
rect 187240 222158 187292 222164
rect 187252 199170 187280 222158
rect 187240 199164 187292 199170
rect 187240 199106 187292 199112
rect 187146 198520 187202 198529
rect 187146 198455 187202 198464
rect 187344 198393 187372 259422
rect 187424 218068 187476 218074
rect 187424 218010 187476 218016
rect 187436 199102 187464 218010
rect 187620 205737 187648 280162
rect 188344 262268 188396 262274
rect 188344 262210 188396 262216
rect 187606 205728 187662 205737
rect 187516 205692 187568 205698
rect 187606 205663 187662 205672
rect 187516 205634 187568 205640
rect 187424 199096 187476 199102
rect 187424 199038 187476 199044
rect 187528 199034 187556 205634
rect 188252 202904 188304 202910
rect 188252 202846 188304 202852
rect 187976 201544 188028 201550
rect 187976 201486 188028 201492
rect 187988 199306 188016 201486
rect 187976 199300 188028 199306
rect 187976 199242 188028 199248
rect 187516 199028 187568 199034
rect 187516 198970 187568 198976
rect 188264 198966 188292 202846
rect 188252 198960 188304 198966
rect 188252 198902 188304 198908
rect 187330 198384 187386 198393
rect 187330 198319 187386 198328
rect 188356 197946 188384 262210
rect 188436 256760 188488 256766
rect 188436 256702 188488 256708
rect 188448 198082 188476 256702
rect 188528 231872 188580 231878
rect 188528 231814 188580 231820
rect 188540 199442 188568 231814
rect 188620 227860 188672 227866
rect 188620 227802 188672 227808
rect 188528 199436 188580 199442
rect 188528 199378 188580 199384
rect 188632 198150 188660 227802
rect 188712 223644 188764 223650
rect 188712 223586 188764 223592
rect 188724 198286 188752 223586
rect 188896 221536 188948 221542
rect 188896 221478 188948 221484
rect 188804 221468 188856 221474
rect 188804 221410 188856 221416
rect 188712 198280 188764 198286
rect 188712 198222 188764 198228
rect 188620 198144 188672 198150
rect 188620 198086 188672 198092
rect 188436 198076 188488 198082
rect 188436 198018 188488 198024
rect 188344 197940 188396 197946
rect 188344 197882 188396 197888
rect 188816 197878 188844 221410
rect 188804 197872 188856 197878
rect 188804 197814 188856 197820
rect 188908 197810 188936 221478
rect 188988 219496 189040 219502
rect 188988 219438 189040 219444
rect 189000 198354 189028 219438
rect 189078 219328 189134 219337
rect 189078 219263 189134 219272
rect 189092 218210 189120 219263
rect 189080 218204 189132 218210
rect 189080 218146 189132 218152
rect 189078 216336 189134 216345
rect 189078 216271 189134 216280
rect 189092 215354 189120 216271
rect 189080 215348 189132 215354
rect 189080 215290 189132 215296
rect 189736 202842 189764 285398
rect 189908 284844 189960 284850
rect 189908 284786 189960 284792
rect 189816 274712 189868 274718
rect 189816 274654 189868 274660
rect 189724 202836 189776 202842
rect 189724 202778 189776 202784
rect 188988 198348 189040 198354
rect 188988 198290 189040 198296
rect 188896 197804 188948 197810
rect 188896 197746 188948 197752
rect 189828 196654 189856 274654
rect 189920 230450 189948 284786
rect 189998 279168 190054 279177
rect 189998 279103 190054 279112
rect 190012 278798 190040 279103
rect 190000 278792 190052 278798
rect 190000 278734 190052 278740
rect 190000 248464 190052 248470
rect 190000 248406 190052 248412
rect 189908 230444 189960 230450
rect 189908 230386 189960 230392
rect 189906 217696 189962 217705
rect 189906 217631 189962 217640
rect 189920 200122 189948 217631
rect 189908 200116 189960 200122
rect 189908 200058 189960 200064
rect 190012 196790 190040 248406
rect 190090 214840 190146 214849
rect 190090 214775 190146 214784
rect 190104 213994 190132 214775
rect 190092 213988 190144 213994
rect 190092 213930 190144 213936
rect 190274 213616 190330 213625
rect 190274 213551 190330 213560
rect 190288 213246 190316 213551
rect 190276 213240 190328 213246
rect 190276 213182 190328 213188
rect 190000 196784 190052 196790
rect 190000 196726 190052 196732
rect 189816 196648 189868 196654
rect 189816 196590 189868 196596
rect 186964 196580 187016 196586
rect 186964 196522 187016 196528
rect 189080 196036 189132 196042
rect 189080 195978 189132 195984
rect 189092 195906 189120 195978
rect 189080 195900 189132 195906
rect 189080 195842 189132 195848
rect 155960 195560 156012 195566
rect 155960 195502 156012 195508
rect 146024 195220 146076 195226
rect 146024 195162 146076 195168
rect 81072 191820 81124 191826
rect 81072 191762 81124 191768
rect 78588 186312 78640 186318
rect 78588 186254 78640 186260
rect 74448 184884 74500 184890
rect 74448 184826 74500 184832
rect 66168 183524 66220 183530
rect 66168 183466 66220 183472
rect 49424 182844 49476 182850
rect 49424 182786 49476 182792
rect 88064 182232 88116 182238
rect 88064 182174 88116 182180
rect 49332 182164 49384 182170
rect 49332 182106 49384 182112
rect 88076 177886 88104 182174
rect 191116 179586 191144 700402
rect 192484 465996 192536 466002
rect 192484 465938 192536 465944
rect 191288 465044 191340 465050
rect 191288 464986 191340 464992
rect 191196 433424 191248 433430
rect 191196 433366 191248 433372
rect 191208 379409 191236 433366
rect 191300 413982 191328 464986
rect 191472 464296 191524 464302
rect 191472 464238 191524 464244
rect 191380 464228 191432 464234
rect 191380 464170 191432 464176
rect 191392 426426 191420 464170
rect 191380 426420 191432 426426
rect 191380 426362 191432 426368
rect 191380 423700 191432 423706
rect 191380 423642 191432 423648
rect 191288 413976 191340 413982
rect 191288 413918 191340 413924
rect 191288 389292 191340 389298
rect 191288 389234 191340 389240
rect 191194 379400 191250 379409
rect 191194 379335 191250 379344
rect 191300 379302 191328 389234
rect 191288 379296 191340 379302
rect 191288 379238 191340 379244
rect 191392 377738 191420 423642
rect 191484 422278 191512 464238
rect 191472 422272 191524 422278
rect 191472 422214 191524 422220
rect 191472 419552 191524 419558
rect 191472 419494 191524 419500
rect 191484 377874 191512 419494
rect 191564 415472 191616 415478
rect 191564 415414 191616 415420
rect 191576 377942 191604 415414
rect 191564 377936 191616 377942
rect 191564 377878 191616 377884
rect 191472 377868 191524 377874
rect 191472 377810 191524 377816
rect 191380 377732 191432 377738
rect 191380 377674 191432 377680
rect 191196 340196 191248 340202
rect 191196 340138 191248 340144
rect 191104 179580 191156 179586
rect 191104 179522 191156 179528
rect 88064 177880 88116 177886
rect 88064 177822 88116 177828
rect 191208 177449 191236 340138
rect 192496 298110 192524 465938
rect 192668 465792 192720 465798
rect 192668 465734 192720 465740
rect 192576 465656 192628 465662
rect 192576 465598 192628 465604
rect 192588 303550 192616 465598
rect 192680 405686 192708 465734
rect 195242 465624 195298 465633
rect 195242 465559 195298 465568
rect 193864 465452 193916 465458
rect 193864 465394 193916 465400
rect 192668 405680 192720 405686
rect 192668 405622 192720 405628
rect 192852 403028 192904 403034
rect 192852 402970 192904 402976
rect 192668 398880 192720 398886
rect 192668 398822 192720 398828
rect 192680 309058 192708 398822
rect 192760 394732 192812 394738
rect 192760 394674 192812 394680
rect 192772 322930 192800 394674
rect 192864 377602 192892 402970
rect 192852 377596 192904 377602
rect 192852 377538 192904 377544
rect 193876 347682 193904 465394
rect 193956 427848 194008 427854
rect 193956 427790 194008 427796
rect 193968 377806 193996 427790
rect 194048 398880 194100 398886
rect 194048 398822 194100 398828
rect 194060 379438 194088 398822
rect 194140 394732 194192 394738
rect 194140 394674 194192 394680
rect 194048 379432 194100 379438
rect 194048 379374 194100 379380
rect 194152 379166 194180 394674
rect 194140 379160 194192 379166
rect 194140 379102 194192 379108
rect 193956 377800 194008 377806
rect 193956 377742 194008 377748
rect 193864 347676 193916 347682
rect 193864 347618 193916 347624
rect 192760 322924 192812 322930
rect 192760 322866 192812 322872
rect 192668 309052 192720 309058
rect 192668 308994 192720 309000
rect 192576 303544 192628 303550
rect 192576 303486 192628 303492
rect 195256 300762 195284 465559
rect 198096 465384 198148 465390
rect 198096 465326 198148 465332
rect 198004 465316 198056 465322
rect 198004 465258 198056 465264
rect 196624 464364 196676 464370
rect 196624 464306 196676 464312
rect 195336 458244 195388 458250
rect 195336 458186 195388 458192
rect 195244 300756 195296 300762
rect 195244 300698 195296 300704
rect 192484 298104 192536 298110
rect 192484 298046 192536 298052
rect 195348 295322 195376 458186
rect 195612 407176 195664 407182
rect 195612 407118 195664 407124
rect 195428 397520 195480 397526
rect 195428 397462 195480 397468
rect 195440 313206 195468 397462
rect 195520 396092 195572 396098
rect 195520 396034 195572 396040
rect 195532 318782 195560 396034
rect 195624 377534 195652 407118
rect 195612 377528 195664 377534
rect 195612 377470 195664 377476
rect 195520 318776 195572 318782
rect 195520 318718 195572 318724
rect 195428 313200 195480 313206
rect 195428 313142 195480 313148
rect 196636 310418 196664 464306
rect 196808 420980 196860 420986
rect 196808 420922 196860 420928
rect 196716 393372 196768 393378
rect 196716 393314 196768 393320
rect 196728 328370 196756 393314
rect 196820 379506 196848 420922
rect 196900 415540 196952 415546
rect 196900 415482 196952 415488
rect 196808 379500 196860 379506
rect 196808 379442 196860 379448
rect 196912 377330 196940 415482
rect 196992 411324 197044 411330
rect 196992 411266 197044 411272
rect 197004 377398 197032 411266
rect 196992 377392 197044 377398
rect 196992 377334 197044 377340
rect 196900 377324 196952 377330
rect 196900 377266 196952 377272
rect 198016 335238 198044 465258
rect 198108 339454 198136 465326
rect 198188 437572 198240 437578
rect 198188 437514 198240 437520
rect 198200 378622 198228 437514
rect 198280 429208 198332 429214
rect 198280 429150 198332 429156
rect 198292 378690 198320 429150
rect 198372 425128 198424 425134
rect 198372 425070 198424 425076
rect 198384 378758 198412 425070
rect 198372 378752 198424 378758
rect 198372 378694 198424 378700
rect 198280 378684 198332 378690
rect 198280 378626 198332 378632
rect 198188 378616 198240 378622
rect 198188 378558 198240 378564
rect 198096 339448 198148 339454
rect 198096 339390 198148 339396
rect 198004 335232 198056 335238
rect 198004 335174 198056 335180
rect 196716 328364 196768 328370
rect 196716 328306 196768 328312
rect 196624 310412 196676 310418
rect 196624 310354 196676 310360
rect 195336 295316 195388 295322
rect 195336 295258 195388 295264
rect 192484 286612 192536 286618
rect 192484 286554 192536 286560
rect 191472 286000 191524 286006
rect 191472 285942 191524 285948
rect 191288 285660 191340 285666
rect 191288 285602 191340 285608
rect 191300 212498 191328 285602
rect 191380 253972 191432 253978
rect 191380 253914 191432 253920
rect 191288 212492 191340 212498
rect 191288 212434 191340 212440
rect 191288 208412 191340 208418
rect 191288 208354 191340 208360
rect 191300 197130 191328 208354
rect 191288 197124 191340 197130
rect 191288 197066 191340 197072
rect 191392 196722 191420 253914
rect 191484 238746 191512 285942
rect 191564 240168 191616 240174
rect 191564 240110 191616 240116
rect 191472 238740 191524 238746
rect 191472 238682 191524 238688
rect 191472 215348 191524 215354
rect 191472 215290 191524 215296
rect 191484 205630 191512 215290
rect 191472 205624 191524 205630
rect 191472 205566 191524 205572
rect 191472 202972 191524 202978
rect 191472 202914 191524 202920
rect 191484 197198 191512 202914
rect 191472 197192 191524 197198
rect 191472 197134 191524 197140
rect 191576 196858 191604 240110
rect 191656 213988 191708 213994
rect 191656 213930 191708 213936
rect 191668 209778 191696 213930
rect 191656 209772 191708 209778
rect 191656 209714 191708 209720
rect 191564 196852 191616 196858
rect 191564 196794 191616 196800
rect 191380 196716 191432 196722
rect 191380 196658 191432 196664
rect 192496 184822 192524 286554
rect 192576 286544 192628 286550
rect 192576 286486 192628 286492
rect 192588 190398 192616 286486
rect 194048 286068 194100 286074
rect 194048 286010 194100 286016
rect 192760 285932 192812 285938
rect 192760 285874 192812 285880
rect 192668 280288 192720 280294
rect 192668 280230 192720 280236
rect 192680 195226 192708 280230
rect 192772 234598 192800 285874
rect 193864 285320 193916 285326
rect 193864 285262 193916 285268
rect 192760 234592 192812 234598
rect 192760 234534 192812 234540
rect 192760 218136 192812 218142
rect 192760 218078 192812 218084
rect 192772 197266 192800 218078
rect 193876 208350 193904 285262
rect 193956 244316 194008 244322
rect 193956 244258 194008 244264
rect 193864 208344 193916 208350
rect 193864 208286 193916 208292
rect 192760 197260 192812 197266
rect 192760 197202 192812 197208
rect 193968 195838 193996 244258
rect 194060 242894 194088 286010
rect 195244 285592 195296 285598
rect 195244 285534 195296 285540
rect 194048 242888 194100 242894
rect 194048 242830 194100 242836
rect 194048 222284 194100 222290
rect 194048 222226 194100 222232
rect 194060 197334 194088 222226
rect 195256 216646 195284 285534
rect 198096 285524 198148 285530
rect 198096 285466 198148 285472
rect 198004 267776 198056 267782
rect 198004 267718 198056 267724
rect 196624 259548 196676 259554
rect 196624 259490 196676 259496
rect 195336 251252 195388 251258
rect 195336 251194 195388 251200
rect 195244 216640 195296 216646
rect 195244 216582 195296 216588
rect 194048 197328 194100 197334
rect 194048 197270 194100 197276
rect 193956 195832 194008 195838
rect 193956 195774 194008 195780
rect 195348 195498 195376 251194
rect 195428 249824 195480 249830
rect 195428 249766 195480 249772
rect 195440 195634 195468 249766
rect 195520 247104 195572 247110
rect 195520 247046 195572 247052
rect 195532 195770 195560 247046
rect 195612 236020 195664 236026
rect 195612 235962 195664 235968
rect 195624 196926 195652 235962
rect 195612 196920 195664 196926
rect 195612 196862 195664 196868
rect 195520 195764 195572 195770
rect 195520 195706 195572 195712
rect 195428 195628 195480 195634
rect 195428 195570 195480 195576
rect 195336 195492 195388 195498
rect 195336 195434 195388 195440
rect 196636 195362 196664 259490
rect 196716 254040 196768 254046
rect 196716 253982 196768 253988
rect 196728 195430 196756 253982
rect 196716 195424 196768 195430
rect 196716 195366 196768 195372
rect 196624 195356 196676 195362
rect 196624 195298 196676 195304
rect 198016 195294 198044 267718
rect 198108 222154 198136 285466
rect 215944 278792 215996 278798
rect 215944 278734 215996 278740
rect 198096 222148 198148 222154
rect 198096 222090 198148 222096
rect 198096 218204 198148 218210
rect 198096 218146 198148 218152
rect 198004 195288 198056 195294
rect 198004 195230 198056 195236
rect 192668 195220 192720 195226
rect 192668 195162 192720 195168
rect 198108 194478 198136 218146
rect 198096 194472 198148 194478
rect 198096 194414 198148 194420
rect 192576 190392 192628 190398
rect 192576 190334 192628 190340
rect 192484 184816 192536 184822
rect 192484 184758 192536 184764
rect 215956 182102 215984 278734
rect 215944 182096 215996 182102
rect 215944 182038 215996 182044
rect 218072 180266 218100 703582
rect 218808 703474 218836 703582
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 218992 703474 219020 703520
rect 218808 703446 219020 703474
rect 233884 700528 233936 700534
rect 233884 700470 233936 700476
rect 228364 305040 228416 305046
rect 228364 304982 228416 304988
rect 218060 180260 218112 180266
rect 218060 180202 218112 180208
rect 228376 177750 228404 304982
rect 232502 285832 232558 285841
rect 232502 285767 232558 285776
rect 228456 209840 228508 209846
rect 228456 209782 228508 209788
rect 228468 198762 228496 209782
rect 228456 198756 228508 198762
rect 228456 198698 228508 198704
rect 232516 191758 232544 285767
rect 232596 285728 232648 285734
rect 232596 285670 232648 285676
rect 232608 197334 232636 285670
rect 232596 197328 232648 197334
rect 232596 197270 232648 197276
rect 232504 191752 232556 191758
rect 232504 191694 232556 191700
rect 233896 179858 233924 700470
rect 239404 700460 239456 700466
rect 239404 700402 239456 700408
rect 233976 656940 234028 656946
rect 233976 656882 234028 656888
rect 233884 179852 233936 179858
rect 233884 179794 233936 179800
rect 233988 179217 234016 656882
rect 238024 466064 238076 466070
rect 238024 466006 238076 466012
rect 235264 464908 235316 464914
rect 235264 464850 235316 464856
rect 235276 321570 235304 464850
rect 235356 464568 235408 464574
rect 235356 464510 235408 464516
rect 235368 325582 235396 464510
rect 237470 438152 237526 438161
rect 237470 438087 237526 438096
rect 237378 437608 237434 437617
rect 237484 437578 237512 438087
rect 237378 437543 237434 437552
rect 237472 437572 237524 437578
rect 237392 437510 237420 437543
rect 237472 437514 237524 437520
rect 237380 437504 237432 437510
rect 237380 437446 237432 437452
rect 237470 433664 237526 433673
rect 237470 433599 237526 433608
rect 237380 433424 237432 433430
rect 237378 433392 237380 433401
rect 237432 433392 237434 433401
rect 237484 433362 237512 433599
rect 237378 433327 237434 433336
rect 237472 433356 237524 433362
rect 237472 433298 237524 433304
rect 237380 431928 237432 431934
rect 237380 431870 237432 431876
rect 237392 431361 237420 431870
rect 237378 431352 237434 431361
rect 237378 431287 237434 431296
rect 237378 429312 237434 429321
rect 237378 429247 237434 429256
rect 237392 429214 237420 429247
rect 237380 429208 237432 429214
rect 237380 429150 237432 429156
rect 237378 428496 237434 428505
rect 237378 428431 237434 428440
rect 237392 427854 237420 428431
rect 237380 427848 237432 427854
rect 237380 427790 237432 427796
rect 237380 426420 237432 426426
rect 237380 426362 237432 426368
rect 237392 426329 237420 426362
rect 237378 426320 237434 426329
rect 237378 426255 237434 426264
rect 237378 425232 237434 425241
rect 237378 425167 237434 425176
rect 237392 425134 237420 425167
rect 237380 425128 237432 425134
rect 237380 425070 237432 425076
rect 237378 424008 237434 424017
rect 237378 423943 237434 423952
rect 237392 423706 237420 423943
rect 237380 423700 237432 423706
rect 237380 423642 237432 423648
rect 237380 422272 237432 422278
rect 237380 422214 237432 422220
rect 237392 422113 237420 422214
rect 237378 422104 237434 422113
rect 237378 422039 237434 422048
rect 237378 421016 237434 421025
rect 237378 420951 237380 420960
rect 237432 420951 237434 420960
rect 237380 420922 237432 420928
rect 237378 419656 237434 419665
rect 237378 419591 237434 419600
rect 237392 419558 237420 419591
rect 237380 419552 237432 419558
rect 237380 419494 237432 419500
rect 237470 416120 237526 416129
rect 237470 416055 237526 416064
rect 237378 415576 237434 415585
rect 237484 415546 237512 416055
rect 237378 415511 237434 415520
rect 237472 415540 237524 415546
rect 237392 415478 237420 415511
rect 237472 415482 237524 415488
rect 237380 415472 237432 415478
rect 237380 415414 237432 415420
rect 237380 413976 237432 413982
rect 237380 413918 237432 413924
rect 237392 413817 237420 413918
rect 237378 413808 237434 413817
rect 237378 413743 237434 413752
rect 237378 411768 237434 411777
rect 237378 411703 237434 411712
rect 237392 411330 237420 411703
rect 237380 411324 237432 411330
rect 237380 411266 237432 411272
rect 237378 407416 237434 407425
rect 237378 407351 237434 407360
rect 237392 407182 237420 407351
rect 237380 407176 237432 407182
rect 237380 407118 237432 407124
rect 237380 405680 237432 405686
rect 237380 405622 237432 405628
rect 237392 405113 237420 405622
rect 237378 405104 237434 405113
rect 237378 405039 237434 405048
rect 237378 403336 237434 403345
rect 237378 403271 237434 403280
rect 237392 403034 237420 403271
rect 237380 403028 237432 403034
rect 237380 402970 237432 402976
rect 237380 400172 237432 400178
rect 237380 400114 237432 400120
rect 237392 400081 237420 400114
rect 237378 400072 237434 400081
rect 237378 400007 237434 400016
rect 237378 398984 237434 398993
rect 237378 398919 237434 398928
rect 237392 398886 237420 398919
rect 237380 398880 237432 398886
rect 237380 398822 237432 398828
rect 237380 396024 237432 396030
rect 237378 395992 237380 396001
rect 237432 395992 237434 396001
rect 237378 395927 237434 395936
rect 237378 394768 237434 394777
rect 237378 394703 237380 394712
rect 237432 394703 237434 394712
rect 237380 394674 237432 394680
rect 237380 391944 237432 391950
rect 237378 391912 237380 391921
rect 237432 391912 237434 391921
rect 237378 391847 237434 391856
rect 237470 389736 237526 389745
rect 237470 389671 237526 389680
rect 237378 389328 237434 389337
rect 237484 389298 237512 389671
rect 237378 389263 237434 389272
rect 237472 389292 237524 389298
rect 237392 389230 237420 389263
rect 237472 389234 237524 389240
rect 237380 389224 237432 389230
rect 237380 389166 237432 389172
rect 237380 387796 237432 387802
rect 237380 387738 237432 387744
rect 237392 387433 237420 387738
rect 237378 387424 237434 387433
rect 237378 387359 237434 387368
rect 237378 385384 237434 385393
rect 237378 385319 237434 385328
rect 237392 385082 237420 385319
rect 237470 385112 237526 385121
rect 237380 385076 237432 385082
rect 237470 385047 237526 385056
rect 237380 385018 237432 385024
rect 237380 383648 237432 383654
rect 237380 383590 237432 383596
rect 237392 383081 237420 383590
rect 237378 383072 237434 383081
rect 237378 383007 237434 383016
rect 237378 381032 237434 381041
rect 237378 380967 237434 380976
rect 237392 380934 237420 380967
rect 237380 380928 237432 380934
rect 237380 380870 237432 380876
rect 237378 380080 237434 380089
rect 237378 380015 237434 380024
rect 237392 378826 237420 380015
rect 237380 378820 237432 378826
rect 237380 378762 237432 378768
rect 237484 378146 237512 385047
rect 237472 378140 237524 378146
rect 237472 378082 237524 378088
rect 237380 377460 237432 377466
rect 237380 377402 237432 377408
rect 237392 377369 237420 377402
rect 237378 377360 237434 377369
rect 237378 377295 237434 377304
rect 237380 376712 237432 376718
rect 237378 376680 237380 376689
rect 237432 376680 237434 376689
rect 237378 376615 237434 376624
rect 237380 373992 237432 373998
rect 237380 373934 237432 373940
rect 237392 373425 237420 373934
rect 237378 373416 237434 373425
rect 237378 373351 237434 373360
rect 237380 372564 237432 372570
rect 237380 372506 237432 372512
rect 237392 372337 237420 372506
rect 237378 372328 237434 372337
rect 237378 372263 237434 372272
rect 237472 368484 237524 368490
rect 237472 368426 237524 368432
rect 237380 368416 237432 368422
rect 237378 368384 237380 368393
rect 237432 368384 237434 368393
rect 237378 368319 237434 368328
rect 237484 368121 237512 368426
rect 237470 368112 237526 368121
rect 237470 368047 237526 368056
rect 238036 365537 238064 466006
rect 238208 465248 238260 465254
rect 238208 465190 238260 465196
rect 238116 465180 238168 465186
rect 238116 465122 238168 465128
rect 238128 369753 238156 465122
rect 238220 373969 238248 465190
rect 238392 464500 238444 464506
rect 238392 464442 238444 464448
rect 238300 464432 238352 464438
rect 238300 464374 238352 464380
rect 238312 409465 238340 464374
rect 238404 418169 238432 464442
rect 238484 463072 238536 463078
rect 238484 463014 238536 463020
rect 238496 435849 238524 463014
rect 238576 463004 238628 463010
rect 238576 462946 238628 462952
rect 238588 440201 238616 462946
rect 238574 440192 238630 440201
rect 238574 440127 238630 440136
rect 239312 436620 239364 436626
rect 239312 436562 239364 436568
rect 238482 435840 238538 435849
rect 238482 435775 238538 435784
rect 238390 418160 238446 418169
rect 238390 418095 238446 418104
rect 238390 411360 238446 411369
rect 238390 411295 238446 411304
rect 238298 409456 238354 409465
rect 238298 409391 238354 409400
rect 238298 406464 238354 406473
rect 238298 406399 238354 406408
rect 238312 378010 238340 406399
rect 238404 379030 238432 411295
rect 238482 402112 238538 402121
rect 238482 402047 238538 402056
rect 238392 379024 238444 379030
rect 238392 378966 238444 378972
rect 238496 378078 238524 402047
rect 238574 397624 238630 397633
rect 238574 397559 238630 397568
rect 238588 378962 238616 397559
rect 238666 393408 238722 393417
rect 238666 393343 238722 393352
rect 238576 378956 238628 378962
rect 238576 378898 238628 378904
rect 238680 378894 238708 393343
rect 238668 378888 238720 378894
rect 238668 378830 238720 378836
rect 238484 378072 238536 378078
rect 238484 378014 238536 378020
rect 238300 378004 238352 378010
rect 238300 377946 238352 377952
rect 238300 376032 238352 376038
rect 238300 375974 238352 375980
rect 238206 373960 238262 373969
rect 238206 373895 238262 373904
rect 238114 369744 238170 369753
rect 238114 369679 238170 369688
rect 238022 365528 238078 365537
rect 238022 365463 238078 365472
rect 237472 364336 237524 364342
rect 237472 364278 237524 364284
rect 237380 364268 237432 364274
rect 237380 364210 237432 364216
rect 237392 364177 237420 364210
rect 237378 364168 237434 364177
rect 237378 364103 237434 364112
rect 237484 363769 237512 364278
rect 237470 363760 237526 363769
rect 237470 363695 237526 363704
rect 237380 361548 237432 361554
rect 237380 361490 237432 361496
rect 237392 361185 237420 361490
rect 237378 361176 237434 361185
rect 237378 361111 237434 361120
rect 237380 360188 237432 360194
rect 237380 360130 237432 360136
rect 237392 359961 237420 360130
rect 237378 359952 237434 359961
rect 237378 359887 237434 359896
rect 237380 358760 237432 358766
rect 237378 358728 237380 358737
rect 237432 358728 237434 358737
rect 237378 358663 237434 358672
rect 237380 356040 237432 356046
rect 237380 355982 237432 355988
rect 237392 355881 237420 355982
rect 237378 355872 237434 355881
rect 237378 355807 237434 355816
rect 237380 354680 237432 354686
rect 237378 354648 237380 354657
rect 237432 354648 237434 354657
rect 237378 354583 237434 354592
rect 237380 351892 237432 351898
rect 237380 351834 237432 351840
rect 237392 351529 237420 351834
rect 237378 351520 237434 351529
rect 237378 351455 237434 351464
rect 237380 350532 237432 350538
rect 237380 350474 237432 350480
rect 237392 350305 237420 350474
rect 237378 350296 237434 350305
rect 237378 350231 237434 350240
rect 237472 347744 237524 347750
rect 237472 347686 237524 347692
rect 237380 347676 237432 347682
rect 237380 347618 237432 347624
rect 237392 347585 237420 347618
rect 237378 347576 237434 347585
rect 237378 347511 237434 347520
rect 237484 347041 237512 347686
rect 238024 347064 238076 347070
rect 237470 347032 237526 347041
rect 238024 347006 238076 347012
rect 237470 346967 237526 346976
rect 237380 346384 237432 346390
rect 237380 346326 237432 346332
rect 237392 346225 237420 346326
rect 237378 346216 237434 346225
rect 237378 346151 237434 346160
rect 237380 343596 237432 343602
rect 237380 343538 237432 343544
rect 237392 343505 237420 343538
rect 237378 343496 237434 343505
rect 237378 343431 237434 343440
rect 237472 342236 237524 342242
rect 237472 342178 237524 342184
rect 237380 342168 237432 342174
rect 237378 342136 237380 342145
rect 237432 342136 237434 342145
rect 237378 342071 237434 342080
rect 237484 341873 237512 342178
rect 237470 341864 237526 341873
rect 237470 341799 237526 341808
rect 237380 339448 237432 339454
rect 237380 339390 237432 339396
rect 237392 339153 237420 339390
rect 237378 339144 237434 339153
rect 237378 339079 237434 339088
rect 237472 338088 237524 338094
rect 237472 338030 237524 338036
rect 237380 338020 237432 338026
rect 237380 337962 237432 337968
rect 237392 337929 237420 337962
rect 237378 337920 237434 337929
rect 237378 337855 237434 337864
rect 237484 337385 237512 338030
rect 237470 337376 237526 337385
rect 237470 337311 237526 337320
rect 237380 336728 237432 336734
rect 237380 336670 237432 336676
rect 237392 336569 237420 336670
rect 237378 336560 237434 336569
rect 237378 336495 237434 336504
rect 237380 335300 237432 335306
rect 237380 335242 237432 335248
rect 237392 335209 237420 335242
rect 237472 335232 237524 335238
rect 237378 335200 237434 335209
rect 237472 335174 237524 335180
rect 237378 335135 237434 335144
rect 237484 334801 237512 335174
rect 237470 334792 237526 334801
rect 237470 334727 237526 334736
rect 237380 333940 237432 333946
rect 237380 333882 237432 333888
rect 237392 333849 237420 333882
rect 237378 333840 237434 333849
rect 237378 333775 237434 333784
rect 237380 332580 237432 332586
rect 237380 332522 237432 332528
rect 237392 332489 237420 332522
rect 237472 332512 237524 332518
rect 237378 332480 237434 332489
rect 237472 332454 237524 332460
rect 237378 332415 237434 332424
rect 237484 332217 237512 332454
rect 237470 332208 237526 332217
rect 237470 332143 237526 332152
rect 237380 331220 237432 331226
rect 237380 331162 237432 331168
rect 237392 330993 237420 331162
rect 237378 330984 237434 330993
rect 237378 330919 237434 330928
rect 237380 329792 237432 329798
rect 237380 329734 237432 329740
rect 237392 329497 237420 329734
rect 237378 329488 237434 329497
rect 237378 329423 237434 329432
rect 237380 328432 237432 328438
rect 237380 328374 237432 328380
rect 237392 328273 237420 328374
rect 237472 328364 237524 328370
rect 237472 328306 237524 328312
rect 237378 328264 237434 328273
rect 237378 328199 237434 328208
rect 237484 327729 237512 328306
rect 237470 327720 237526 327729
rect 237470 327655 237526 327664
rect 237380 327072 237432 327078
rect 237380 327014 237432 327020
rect 237392 326913 237420 327014
rect 237378 326904 237434 326913
rect 237378 326839 237434 326848
rect 237380 325644 237432 325650
rect 237380 325586 237432 325592
rect 235356 325576 235408 325582
rect 235356 325518 235408 325524
rect 237392 325145 237420 325586
rect 237472 325576 237524 325582
rect 237470 325544 237472 325553
rect 237524 325544 237526 325553
rect 237470 325479 237526 325488
rect 237378 325136 237434 325145
rect 237378 325071 237434 325080
rect 237380 324284 237432 324290
rect 237380 324226 237432 324232
rect 237392 324193 237420 324226
rect 237378 324184 237434 324193
rect 237378 324119 237434 324128
rect 237380 322924 237432 322930
rect 237380 322866 237432 322872
rect 237392 322833 237420 322866
rect 237378 322824 237434 322833
rect 237378 322759 237434 322768
rect 235264 321564 235316 321570
rect 235264 321506 235316 321512
rect 237380 321564 237432 321570
rect 237380 321506 237432 321512
rect 237392 321473 237420 321506
rect 237378 321464 237434 321473
rect 237378 321399 237434 321408
rect 237472 320136 237524 320142
rect 237378 320104 237434 320113
rect 237472 320078 237524 320084
rect 237378 320039 237380 320048
rect 237432 320039 237434 320048
rect 237380 320010 237432 320016
rect 237484 319841 237512 320078
rect 237470 319832 237526 319841
rect 237470 319767 237526 319776
rect 237380 318776 237432 318782
rect 237380 318718 237432 318724
rect 237392 318617 237420 318718
rect 237378 318608 237434 318617
rect 237378 318543 237434 318552
rect 238036 318073 238064 347006
rect 238312 322425 238340 375974
rect 238298 322416 238354 322425
rect 238298 322351 238354 322360
rect 238022 318064 238078 318073
rect 238022 317999 238078 318008
rect 237380 317416 237432 317422
rect 237380 317358 237432 317364
rect 237392 317257 237420 317358
rect 237378 317248 237434 317257
rect 237378 317183 237434 317192
rect 237380 315988 237432 315994
rect 237380 315930 237432 315936
rect 237392 315489 237420 315930
rect 237378 315480 237434 315489
rect 237378 315415 237434 315424
rect 237380 314628 237432 314634
rect 237380 314570 237432 314576
rect 237392 314537 237420 314570
rect 237378 314528 237434 314537
rect 237378 314463 237434 314472
rect 237472 313268 237524 313274
rect 237472 313210 237524 313216
rect 237380 313200 237432 313206
rect 237378 313168 237380 313177
rect 237432 313168 237434 313177
rect 237378 313103 237434 313112
rect 237484 312769 237512 313210
rect 237470 312760 237526 312769
rect 237470 312695 237526 312704
rect 237380 311840 237432 311846
rect 237378 311808 237380 311817
rect 237432 311808 237434 311817
rect 237378 311743 237434 311752
rect 237472 310480 237524 310486
rect 237378 310448 237434 310457
rect 237472 310422 237524 310428
rect 237378 310383 237380 310392
rect 237432 310383 237434 310392
rect 237380 310354 237432 310360
rect 237484 310185 237512 310422
rect 237470 310176 237526 310185
rect 237470 310111 237526 310120
rect 237380 309120 237432 309126
rect 237380 309062 237432 309068
rect 237392 308961 237420 309062
rect 237472 309052 237524 309058
rect 237472 308994 237524 309000
rect 237378 308952 237434 308961
rect 237378 308887 237434 308896
rect 237484 308417 237512 308994
rect 237470 308408 237526 308417
rect 237470 308343 237526 308352
rect 237380 307760 237432 307766
rect 237380 307702 237432 307708
rect 237392 307601 237420 307702
rect 237378 307592 237434 307601
rect 237378 307527 237434 307536
rect 237380 306332 237432 306338
rect 237380 306274 237432 306280
rect 237392 306241 237420 306274
rect 237472 306264 237524 306270
rect 237378 306232 237434 306241
rect 237472 306206 237524 306212
rect 237378 306167 237434 306176
rect 237484 305833 237512 306206
rect 237470 305824 237526 305833
rect 237470 305759 237526 305768
rect 237380 304972 237432 304978
rect 237380 304914 237432 304920
rect 237392 304881 237420 304914
rect 237378 304872 237434 304881
rect 237378 304807 237434 304816
rect 237380 303612 237432 303618
rect 237380 303554 237432 303560
rect 237392 303521 237420 303554
rect 237472 303544 237524 303550
rect 237378 303512 237434 303521
rect 237472 303486 237524 303492
rect 237378 303447 237434 303456
rect 237484 303113 237512 303486
rect 237470 303104 237526 303113
rect 237470 303039 237526 303048
rect 237380 302184 237432 302190
rect 237378 302152 237380 302161
rect 237432 302152 237434 302161
rect 237378 302087 237434 302096
rect 237380 300824 237432 300830
rect 237378 300792 237380 300801
rect 237432 300792 237434 300801
rect 237378 300727 237434 300736
rect 237472 300756 237524 300762
rect 237472 300698 237524 300704
rect 237484 300529 237512 300698
rect 237470 300520 237526 300529
rect 237470 300455 237526 300464
rect 237472 299464 237524 299470
rect 237472 299406 237524 299412
rect 237380 299396 237432 299402
rect 237380 299338 237432 299344
rect 237392 299305 237420 299338
rect 237378 299296 237434 299305
rect 237378 299231 237434 299240
rect 237484 298761 237512 299406
rect 237470 298752 237526 298761
rect 237470 298687 237526 298696
rect 237380 298104 237432 298110
rect 237380 298046 237432 298052
rect 237392 297945 237420 298046
rect 237378 297936 237434 297945
rect 237378 297871 237434 297880
rect 237380 296676 237432 296682
rect 237380 296618 237432 296624
rect 237392 296585 237420 296618
rect 237472 296608 237524 296614
rect 237378 296576 237434 296585
rect 237472 296550 237524 296556
rect 237378 296511 237434 296520
rect 237484 296177 237512 296550
rect 237470 296168 237526 296177
rect 237470 296103 237526 296112
rect 237380 295316 237432 295322
rect 237380 295258 237432 295264
rect 237392 295225 237420 295258
rect 237378 295216 237434 295225
rect 237378 295151 237434 295160
rect 237380 293956 237432 293962
rect 237380 293898 237432 293904
rect 237392 293865 237420 293898
rect 237378 293856 237434 293865
rect 237378 293791 237434 293800
rect 237378 292768 237434 292777
rect 237378 292703 237434 292712
rect 237392 292670 237420 292703
rect 237380 292664 237432 292670
rect 237380 292606 237432 292612
rect 236644 292596 236696 292602
rect 236644 292538 236696 292544
rect 235264 291236 235316 291242
rect 235264 291178 235316 291184
rect 235172 220856 235224 220862
rect 235172 220798 235224 220804
rect 234988 212560 235040 212566
rect 234988 212502 235040 212508
rect 235000 199753 235028 212502
rect 234986 199744 235042 199753
rect 234986 199679 235042 199688
rect 235184 199617 235212 220798
rect 235170 199608 235226 199617
rect 235170 199543 235226 199552
rect 235276 195566 235304 291178
rect 235356 288516 235408 288522
rect 235356 288458 235408 288464
rect 235368 195702 235396 288458
rect 235448 288448 235500 288454
rect 235448 288390 235500 288396
rect 235460 197169 235488 288390
rect 235540 285796 235592 285802
rect 235540 285738 235592 285744
rect 235446 197160 235502 197169
rect 235446 197095 235502 197104
rect 235552 196994 235580 285738
rect 235632 285728 235684 285734
rect 235632 285670 235684 285676
rect 235644 199374 235672 285670
rect 235816 283008 235868 283014
rect 235816 282950 235868 282956
rect 235724 282940 235776 282946
rect 235724 282882 235776 282888
rect 235632 199368 235684 199374
rect 235632 199310 235684 199316
rect 235736 197062 235764 282882
rect 235828 198218 235856 282950
rect 235908 256828 235960 256834
rect 235908 256770 235960 256776
rect 235920 198490 235948 256770
rect 235908 198484 235960 198490
rect 235908 198426 235960 198432
rect 235816 198212 235868 198218
rect 235816 198154 235868 198160
rect 235724 197056 235776 197062
rect 235724 196998 235776 197004
rect 235540 196988 235592 196994
rect 235540 196930 235592 196936
rect 235356 195696 235408 195702
rect 235356 195638 235408 195644
rect 235264 195560 235316 195566
rect 235264 195502 235316 195508
rect 233974 179208 234030 179217
rect 233974 179143 234030 179152
rect 236656 178974 236684 292538
rect 237378 291408 237434 291417
rect 237378 291343 237434 291352
rect 237392 291242 237420 291343
rect 237380 291236 237432 291242
rect 237380 291178 237432 291184
rect 237378 290048 237434 290057
rect 237378 289983 237434 289992
rect 237392 289882 237420 289983
rect 237380 289876 237432 289882
rect 237380 289818 237432 289824
rect 237470 288688 237526 288697
rect 237470 288623 237526 288632
rect 237378 288552 237434 288561
rect 237484 288522 237512 288623
rect 237378 288487 237434 288496
rect 237472 288516 237524 288522
rect 237392 288454 237420 288487
rect 237472 288458 237524 288464
rect 237380 288448 237432 288454
rect 237380 288390 237432 288396
rect 237378 287192 237434 287201
rect 237378 287127 237434 287136
rect 237392 287094 237420 287127
rect 237380 287088 237432 287094
rect 237380 287030 237432 287036
rect 237378 286104 237434 286113
rect 237378 286039 237434 286048
rect 237392 285734 237420 286039
rect 238116 285932 238168 285938
rect 238116 285874 238168 285880
rect 237470 285832 237526 285841
rect 237470 285767 237472 285776
rect 237524 285767 237526 285776
rect 237472 285738 237524 285744
rect 237380 285728 237432 285734
rect 237380 285670 237432 285676
rect 237840 285388 237892 285394
rect 237840 285330 237892 285336
rect 237380 284912 237432 284918
rect 237378 284880 237380 284889
rect 237432 284880 237434 284889
rect 237378 284815 237434 284824
rect 237378 283520 237434 283529
rect 237378 283455 237434 283464
rect 237392 283014 237420 283455
rect 237380 283008 237432 283014
rect 237380 282950 237432 282956
rect 237470 282976 237526 282985
rect 237470 282911 237472 282920
rect 237524 282911 237526 282920
rect 237472 282882 237524 282888
rect 237380 282872 237432 282878
rect 237378 282840 237380 282849
rect 237432 282840 237434 282849
rect 237378 282775 237434 282784
rect 237378 280800 237434 280809
rect 237378 280735 237434 280744
rect 237392 280294 237420 280735
rect 237470 280392 237526 280401
rect 237470 280327 237526 280336
rect 237380 280288 237432 280294
rect 237380 280230 237432 280236
rect 237484 280226 237512 280327
rect 237472 280220 237524 280226
rect 237472 280162 237524 280168
rect 237380 280152 237432 280158
rect 237380 280094 237432 280100
rect 237392 279857 237420 280094
rect 237378 279848 237434 279857
rect 237378 279783 237434 279792
rect 237380 277364 237432 277370
rect 237380 277306 237432 277312
rect 237392 277273 237420 277306
rect 237378 277264 237434 277273
rect 237378 277199 237434 277208
rect 237470 275088 237526 275097
rect 237470 275023 237526 275032
rect 237484 274718 237512 275023
rect 237472 274712 237524 274718
rect 237472 274654 237524 274660
rect 237380 274644 237432 274650
rect 237380 274586 237432 274592
rect 237392 274553 237420 274586
rect 237378 274544 237434 274553
rect 237378 274479 237434 274488
rect 237380 271856 237432 271862
rect 237378 271824 237380 271833
rect 237432 271824 237434 271833
rect 237378 271759 237434 271768
rect 237852 269793 237880 285330
rect 238024 284980 238076 284986
rect 238024 284922 238076 284928
rect 237838 269784 237894 269793
rect 237838 269719 237894 269728
rect 237378 267880 237434 267889
rect 237378 267815 237434 267824
rect 237392 267782 237420 267815
rect 237380 267776 237432 267782
rect 237380 267718 237432 267724
rect 237378 262440 237434 262449
rect 237378 262375 237434 262384
rect 237392 262274 237420 262375
rect 237380 262268 237432 262274
rect 237380 262210 237432 262216
rect 237472 262200 237524 262206
rect 237472 262142 237524 262148
rect 237378 262032 237434 262041
rect 237378 261967 237434 261976
rect 237392 260914 237420 261967
rect 237484 261905 237512 262142
rect 237470 261896 237526 261905
rect 237470 261831 237526 261840
rect 237380 260908 237432 260914
rect 237380 260850 237432 260856
rect 237378 259720 237434 259729
rect 237378 259655 237434 259664
rect 237392 259554 237420 259655
rect 237470 259584 237526 259593
rect 237380 259548 237432 259554
rect 237470 259519 237526 259528
rect 237380 259490 237432 259496
rect 237484 259486 237512 259519
rect 237472 259480 237524 259486
rect 237472 259422 237524 259428
rect 237380 259412 237432 259418
rect 237380 259354 237432 259360
rect 237392 259185 237420 259354
rect 237378 259176 237434 259185
rect 237378 259111 237434 259120
rect 237378 257136 237434 257145
rect 237378 257071 237434 257080
rect 237392 256766 237420 257071
rect 237470 256864 237526 256873
rect 237470 256799 237472 256808
rect 237524 256799 237526 256808
rect 237472 256770 237524 256776
rect 237380 256760 237432 256766
rect 237380 256702 237432 256708
rect 237470 254552 237526 254561
rect 237470 254487 237526 254496
rect 237378 254144 237434 254153
rect 237378 254079 237434 254088
rect 237392 253978 237420 254079
rect 237484 254046 237512 254487
rect 237472 254040 237524 254046
rect 237472 253982 237524 253988
rect 237380 253972 237432 253978
rect 237380 253914 237432 253920
rect 237378 251832 237434 251841
rect 237378 251767 237434 251776
rect 237392 251258 237420 251767
rect 237380 251252 237432 251258
rect 237380 251194 237432 251200
rect 237378 249928 237434 249937
rect 237378 249863 237434 249872
rect 237392 249830 237420 249863
rect 237380 249824 237432 249830
rect 237380 249766 237432 249772
rect 237378 248568 237434 248577
rect 237378 248503 237434 248512
rect 237392 248470 237420 248503
rect 237380 248464 237432 248470
rect 237380 248406 237432 248412
rect 237380 247104 237432 247110
rect 237378 247072 237380 247081
rect 237432 247072 237434 247081
rect 237378 247007 237434 247016
rect 237378 244488 237434 244497
rect 237378 244423 237434 244432
rect 237392 244322 237420 244423
rect 237380 244316 237432 244322
rect 237380 244258 237432 244264
rect 237380 242888 237432 242894
rect 237378 242856 237380 242865
rect 237432 242856 237434 242865
rect 237378 242791 237434 242800
rect 237378 241632 237434 241641
rect 237378 241567 237434 241576
rect 237392 241534 237420 241567
rect 237380 241528 237432 241534
rect 237380 241470 237432 241476
rect 237378 240408 237434 240417
rect 237378 240343 237434 240352
rect 237392 240174 237420 240343
rect 237380 240168 237432 240174
rect 237380 240110 237432 240116
rect 237380 238740 237432 238746
rect 237380 238682 237432 238688
rect 237392 238649 237420 238682
rect 237378 238640 237434 238649
rect 237378 238575 237434 238584
rect 237378 236056 237434 236065
rect 237378 235991 237380 236000
rect 237432 235991 237434 236000
rect 237380 235962 237432 235968
rect 237380 234592 237432 234598
rect 237380 234534 237432 234540
rect 237392 234297 237420 234534
rect 237378 234288 237434 234297
rect 237378 234223 237434 234232
rect 237378 232520 237434 232529
rect 237378 232455 237434 232464
rect 237392 231878 237420 232455
rect 237380 231872 237432 231878
rect 237380 231814 237432 231820
rect 237380 230444 237432 230450
rect 237380 230386 237432 230392
rect 237392 230217 237420 230386
rect 237378 230208 237434 230217
rect 237378 230143 237434 230152
rect 237470 228168 237526 228177
rect 237470 228103 237526 228112
rect 237484 227866 237512 228103
rect 237472 227860 237524 227866
rect 237472 227802 237524 227808
rect 237380 227792 237432 227798
rect 237378 227760 237380 227769
rect 237432 227760 237434 227769
rect 237378 227695 237434 227704
rect 238036 225865 238064 284922
rect 238128 253881 238156 285874
rect 238208 285864 238260 285870
rect 238208 285806 238260 285812
rect 238114 253872 238170 253881
rect 238114 253807 238170 253816
rect 238114 251424 238170 251433
rect 238114 251359 238170 251368
rect 238022 225856 238078 225865
rect 238022 225791 238078 225800
rect 237378 223680 237434 223689
rect 237378 223615 237380 223624
rect 237432 223615 237434 223624
rect 237380 223586 237432 223592
rect 237470 222864 237526 222873
rect 237470 222799 237526 222808
rect 237378 222320 237434 222329
rect 237378 222255 237380 222264
rect 237432 222255 237434 222264
rect 237380 222226 237432 222232
rect 237484 222222 237512 222799
rect 237472 222216 237524 222222
rect 237472 222158 237524 222164
rect 237380 222148 237432 222154
rect 237380 222090 237432 222096
rect 237392 221513 237420 222090
rect 237470 221640 237526 221649
rect 237470 221575 237526 221584
rect 237378 221504 237434 221513
rect 237378 221439 237434 221448
rect 237484 220862 237512 221575
rect 237472 220856 237524 220862
rect 237472 220798 237524 220804
rect 237378 219600 237434 219609
rect 237378 219535 237434 219544
rect 237392 219502 237420 219535
rect 237380 219496 237432 219502
rect 237380 219438 237432 219444
rect 237470 218512 237526 218521
rect 237470 218447 237526 218456
rect 237380 218136 237432 218142
rect 237378 218104 237380 218113
rect 237432 218104 237434 218113
rect 237484 218074 237512 218447
rect 237378 218039 237434 218048
rect 237472 218068 237524 218074
rect 237472 218010 237524 218016
rect 237380 216640 237432 216646
rect 237380 216582 237432 216588
rect 237392 216481 237420 216582
rect 237378 216472 237434 216481
rect 237378 216407 237434 216416
rect 238022 215384 238078 215393
rect 238022 215319 238078 215328
rect 237378 213480 237434 213489
rect 237378 213415 237434 213424
rect 237392 213246 237420 213415
rect 237380 213240 237432 213246
rect 237380 213182 237432 213188
rect 237470 212800 237526 212809
rect 237470 212735 237526 212744
rect 237484 212566 237512 212735
rect 237472 212560 237524 212566
rect 237472 212502 237524 212508
rect 237380 212492 237432 212498
rect 237380 212434 237432 212440
rect 237392 212401 237420 212434
rect 237378 212392 237434 212401
rect 237378 212327 237434 212336
rect 237470 209944 237526 209953
rect 237470 209879 237526 209888
rect 237484 209846 237512 209879
rect 237472 209840 237524 209846
rect 237472 209782 237524 209788
rect 237380 209772 237432 209778
rect 237380 209714 237432 209720
rect 237392 209681 237420 209714
rect 237378 209672 237434 209681
rect 237378 209607 237434 209616
rect 237378 208448 237434 208457
rect 237378 208383 237380 208392
rect 237432 208383 237434 208392
rect 237380 208354 237432 208360
rect 237472 208344 237524 208350
rect 237470 208312 237472 208321
rect 237524 208312 237526 208321
rect 237470 208247 237526 208256
rect 237930 206136 237986 206145
rect 237930 206071 237986 206080
rect 237470 205864 237526 205873
rect 237470 205799 237526 205808
rect 237484 205698 237512 205799
rect 237472 205692 237524 205698
rect 237472 205634 237524 205640
rect 237380 205624 237432 205630
rect 237378 205592 237380 205601
rect 237432 205592 237434 205601
rect 237378 205527 237434 205536
rect 237378 203552 237434 203561
rect 237378 203487 237434 203496
rect 237392 202978 237420 203487
rect 237470 203008 237526 203017
rect 237380 202972 237432 202978
rect 237470 202943 237526 202952
rect 237380 202914 237432 202920
rect 237484 202910 237512 202943
rect 237472 202904 237524 202910
rect 237472 202846 237524 202852
rect 237380 202836 237432 202842
rect 237380 202778 237432 202784
rect 237392 202609 237420 202778
rect 237378 202600 237434 202609
rect 237378 202535 237434 202544
rect 237380 201544 237432 201550
rect 237378 201512 237380 201521
rect 237432 201512 237434 201521
rect 237378 201447 237434 201456
rect 237470 200152 237526 200161
rect 237380 200116 237432 200122
rect 237470 200087 237526 200096
rect 237380 200058 237432 200064
rect 237392 200025 237420 200058
rect 237378 200016 237434 200025
rect 237378 199951 237434 199960
rect 237484 199578 237512 200087
rect 237472 199572 237524 199578
rect 237472 199514 237524 199520
rect 237944 198830 237972 206071
rect 237932 198824 237984 198830
rect 237932 198766 237984 198772
rect 238036 198558 238064 215319
rect 238024 198552 238076 198558
rect 238024 198494 238076 198500
rect 237380 198008 237432 198014
rect 237378 197976 237380 197985
rect 237432 197976 237434 197985
rect 237378 197911 237434 197920
rect 237380 197328 237432 197334
rect 237378 197296 237380 197305
rect 237432 197296 237434 197305
rect 237378 197231 237434 197240
rect 238128 196450 238156 251359
rect 238220 248305 238248 285806
rect 238484 285252 238536 285258
rect 238484 285194 238536 285200
rect 238392 285048 238444 285054
rect 238392 284990 238444 284996
rect 238298 270736 238354 270745
rect 238298 270671 238354 270680
rect 238206 248296 238262 248305
rect 238206 248231 238262 248240
rect 238206 245712 238262 245721
rect 238206 245647 238262 245656
rect 238220 196518 238248 245647
rect 238312 221542 238340 270671
rect 238404 245585 238432 284990
rect 238496 267209 238524 285194
rect 238668 285184 238720 285190
rect 238668 285126 238720 285132
rect 238576 285116 238628 285122
rect 238576 285058 238628 285064
rect 238482 267200 238538 267209
rect 238482 267135 238538 267144
rect 238482 265024 238538 265033
rect 238482 264959 238538 264968
rect 238390 245576 238446 245585
rect 238390 245511 238446 245520
rect 238390 243128 238446 243137
rect 238390 243063 238446 243072
rect 238300 221536 238352 221542
rect 238300 221478 238352 221484
rect 238298 214024 238354 214033
rect 238298 213959 238354 213968
rect 238312 199510 238340 213959
rect 238300 199504 238352 199510
rect 238300 199446 238352 199452
rect 238404 198626 238432 243063
rect 238496 221474 238524 264959
rect 238588 250889 238616 285058
rect 238680 264081 238708 285126
rect 238666 264072 238722 264081
rect 238666 264007 238722 264016
rect 238574 250880 238630 250889
rect 238574 250815 238630 250824
rect 238574 237416 238630 237425
rect 238574 237351 238630 237360
rect 238484 221468 238536 221474
rect 238484 221410 238536 221416
rect 238482 211168 238538 211177
rect 238482 211103 238538 211112
rect 238496 198898 238524 211103
rect 238484 198892 238536 198898
rect 238484 198834 238536 198840
rect 238392 198620 238444 198626
rect 238392 198562 238444 198568
rect 238588 198422 238616 237351
rect 238666 232112 238722 232121
rect 238666 232047 238722 232056
rect 238680 198694 238708 232047
rect 238668 198688 238720 198694
rect 238668 198630 238720 198636
rect 238576 198416 238628 198422
rect 238576 198358 238628 198364
rect 238208 196512 238260 196518
rect 238208 196454 238260 196460
rect 238116 196444 238168 196450
rect 238116 196386 238168 196392
rect 237470 196072 237526 196081
rect 237470 196007 237472 196016
rect 237524 196007 237526 196016
rect 237472 195978 237524 195984
rect 237380 195968 237432 195974
rect 237378 195936 237380 195945
rect 237432 195936 237434 195945
rect 237378 195871 237434 195880
rect 237472 194540 237524 194546
rect 237472 194482 237524 194488
rect 237380 194472 237432 194478
rect 237378 194440 237380 194449
rect 237432 194440 237434 194449
rect 237378 194375 237434 194384
rect 237484 194177 237512 194482
rect 237470 194168 237526 194177
rect 237470 194103 237526 194112
rect 237380 193180 237432 193186
rect 237380 193122 237432 193128
rect 237392 192953 237420 193122
rect 237378 192944 237434 192953
rect 237378 192879 237434 192888
rect 237380 191820 237432 191826
rect 237380 191762 237432 191768
rect 237392 191593 237420 191762
rect 237472 191752 237524 191758
rect 237470 191720 237472 191729
rect 237524 191720 237526 191729
rect 237470 191655 237526 191664
rect 237378 191584 237434 191593
rect 237378 191519 237434 191528
rect 237380 190460 237432 190466
rect 237380 190402 237432 190408
rect 237392 190369 237420 190402
rect 237472 190392 237524 190398
rect 237378 190360 237434 190369
rect 237472 190334 237524 190340
rect 237378 190295 237434 190304
rect 237484 189825 237512 190334
rect 237470 189816 237526 189825
rect 237470 189751 237526 189760
rect 237380 189032 237432 189038
rect 237378 189000 237380 189009
rect 237432 189000 237434 189009
rect 237378 188935 237434 188944
rect 237380 187672 237432 187678
rect 237378 187640 237380 187649
rect 237432 187640 237434 187649
rect 237378 187575 237434 187584
rect 237380 186312 237432 186318
rect 237378 186280 237380 186289
rect 237432 186280 237434 186289
rect 237378 186215 237434 186224
rect 237378 184920 237434 184929
rect 237378 184855 237380 184864
rect 237432 184855 237434 184864
rect 237380 184826 237432 184832
rect 237472 184816 237524 184822
rect 237472 184758 237524 184764
rect 237484 184521 237512 184758
rect 237470 184512 237526 184521
rect 237470 184447 237526 184456
rect 237380 183524 237432 183530
rect 237380 183466 237432 183472
rect 237392 183297 237420 183466
rect 237378 183288 237434 183297
rect 237378 183223 237434 183232
rect 237564 182844 237616 182850
rect 237564 182786 237616 182792
rect 237380 182164 237432 182170
rect 237380 182106 237432 182112
rect 237392 182073 237420 182106
rect 237472 182096 237524 182102
rect 237378 182064 237434 182073
rect 237472 182038 237524 182044
rect 237378 181999 237434 182008
rect 237484 181937 237512 182038
rect 237470 181928 237526 181937
rect 237470 181863 237526 181872
rect 237380 181552 237432 181558
rect 237380 181494 237432 181500
rect 236644 178968 236696 178974
rect 236644 178910 236696 178916
rect 228364 177744 228416 177750
rect 228364 177686 228416 177692
rect 237392 177585 237420 181494
rect 237576 180713 237604 182786
rect 238760 181484 238812 181490
rect 238760 181426 238812 181432
rect 237562 180704 237618 180713
rect 237562 180639 237618 180648
rect 238772 177721 238800 181426
rect 239324 178770 239352 436562
rect 239312 178764 239364 178770
rect 239312 178706 239364 178712
rect 239416 178566 239444 700402
rect 239588 700392 239640 700398
rect 239588 700334 239640 700340
rect 262220 700392 262272 700398
rect 262220 700334 262272 700340
rect 239496 700324 239548 700330
rect 239496 700266 239548 700272
rect 239508 178945 239536 700266
rect 239494 178936 239550 178945
rect 239494 178871 239550 178880
rect 239600 178634 239628 700334
rect 262128 700324 262180 700330
rect 262128 700266 262180 700272
rect 261944 696992 261996 696998
rect 261944 696934 261996 696940
rect 261956 694142 261984 696934
rect 259460 694136 259512 694142
rect 259460 694078 259512 694084
rect 261944 694136 261996 694142
rect 261944 694078 261996 694084
rect 257344 691416 257396 691422
rect 257344 691358 257396 691364
rect 253204 683188 253256 683194
rect 253204 683130 253256 683136
rect 251824 610496 251876 610502
rect 251824 610438 251876 610444
rect 239680 605872 239732 605878
rect 239680 605814 239732 605820
rect 239692 179790 239720 605814
rect 251836 590714 251864 610438
rect 251824 590708 251876 590714
rect 251824 590650 251876 590656
rect 249064 590640 249116 590646
rect 249064 590582 249116 590588
rect 239772 553444 239824 553450
rect 239772 553386 239824 553392
rect 239680 179784 239732 179790
rect 239680 179726 239732 179732
rect 239784 179654 239812 553386
rect 247684 520328 247736 520334
rect 247684 520270 247736 520276
rect 246304 503668 246356 503674
rect 246304 503610 246356 503616
rect 239864 501016 239916 501022
rect 239864 500958 239916 500964
rect 239772 179648 239824 179654
rect 239772 179590 239824 179596
rect 239876 179518 239904 500958
rect 244924 474020 244976 474026
rect 244924 473962 244976 473968
rect 242532 445868 242584 445874
rect 242532 445810 242584 445816
rect 240232 443420 240284 443426
rect 240232 443362 240284 443368
rect 240140 442468 240192 442474
rect 240140 442410 240192 442416
rect 240048 440904 240100 440910
rect 240048 440846 240100 440852
rect 239956 438932 240008 438938
rect 239956 438874 240008 438880
rect 239864 179512 239916 179518
rect 239864 179454 239916 179460
rect 239968 178838 239996 438874
rect 239956 178832 240008 178838
rect 239956 178774 240008 178780
rect 239588 178628 239640 178634
rect 239588 178570 239640 178576
rect 239404 178560 239456 178566
rect 239404 178502 239456 178508
rect 238758 177712 238814 177721
rect 238758 177647 238814 177656
rect 237378 177576 237434 177585
rect 237378 177511 237434 177520
rect 191194 177440 191250 177449
rect 191194 177375 191250 177384
rect 240060 177274 240088 440846
rect 240152 438938 240180 442410
rect 240140 438932 240192 438938
rect 240140 438874 240192 438880
rect 240244 436626 240272 443362
rect 242544 442474 242572 445810
rect 244936 444514 244964 473962
rect 245016 455388 245068 455394
rect 245016 455330 245068 455336
rect 245028 445874 245056 455330
rect 246316 452606 246344 503610
rect 247696 455394 247724 520270
rect 249076 503674 249104 590582
rect 253216 563106 253244 683130
rect 257356 668642 257384 691358
rect 259472 687290 259500 694078
rect 262140 694074 262168 700266
rect 262232 696998 262260 700334
rect 267660 697610 267688 703520
rect 283852 702434 283880 703520
rect 282932 702406 283880 702434
rect 266360 697604 266412 697610
rect 266360 697546 266412 697552
rect 267648 697604 267700 697610
rect 267648 697546 267700 697552
rect 262220 696992 262272 696998
rect 262220 696934 262272 696940
rect 259552 694068 259604 694074
rect 259552 694010 259604 694016
rect 262128 694068 262180 694074
rect 262128 694010 262180 694016
rect 259564 691422 259592 694010
rect 259552 691416 259604 691422
rect 259552 691358 259604 691364
rect 259380 687262 259500 687290
rect 259380 683194 259408 687262
rect 259368 683188 259420 683194
rect 259368 683130 259420 683136
rect 256056 668636 256108 668642
rect 256056 668578 256108 668584
rect 257344 668636 257396 668642
rect 257344 668578 257396 668584
rect 256068 664970 256096 668578
rect 254584 664964 254636 664970
rect 254584 664906 254636 664912
rect 256056 664964 256108 664970
rect 256056 664906 256108 664912
rect 254596 619614 254624 664906
rect 253296 619608 253348 619614
rect 253296 619550 253348 619556
rect 254584 619608 254636 619614
rect 254584 619550 254636 619556
rect 253308 610502 253336 619550
rect 253296 610496 253348 610502
rect 253296 610438 253348 610444
rect 251824 563100 251876 563106
rect 251824 563042 251876 563048
rect 253204 563100 253256 563106
rect 253204 563042 253256 563048
rect 251836 524482 251864 563042
rect 260104 540252 260156 540258
rect 260104 540194 260156 540200
rect 260116 525842 260144 540194
rect 258724 525836 258776 525842
rect 258724 525778 258776 525784
rect 260104 525836 260156 525842
rect 260104 525778 260156 525784
rect 249432 524476 249484 524482
rect 249432 524418 249484 524424
rect 251824 524476 251876 524482
rect 251824 524418 251876 524424
rect 249444 520334 249472 524418
rect 249432 520328 249484 520334
rect 249432 520270 249484 520276
rect 258736 506734 258764 525778
rect 257344 506728 257396 506734
rect 257344 506670 257396 506676
rect 258724 506728 258776 506734
rect 258724 506670 258776 506676
rect 249064 503668 249116 503674
rect 249064 503610 249116 503616
rect 257356 496874 257384 506670
rect 253940 496868 253992 496874
rect 253940 496810 253992 496816
rect 257344 496868 257396 496874
rect 257344 496810 257396 496816
rect 253952 490618 253980 496810
rect 247776 490612 247828 490618
rect 247776 490554 247828 490560
rect 253940 490612 253992 490618
rect 253940 490554 253992 490560
rect 247788 474026 247816 490554
rect 247776 474020 247828 474026
rect 247776 473962 247828 473968
rect 247684 455388 247736 455394
rect 247684 455330 247736 455336
rect 245108 452600 245160 452606
rect 245108 452542 245160 452548
rect 246304 452600 246356 452606
rect 246304 452542 246356 452548
rect 245016 445868 245068 445874
rect 245016 445810 245068 445816
rect 242900 444508 242952 444514
rect 242900 444450 242952 444456
rect 244924 444508 244976 444514
rect 244924 444450 244976 444456
rect 242532 442468 242584 442474
rect 242532 442410 242584 442416
rect 242912 442338 242940 444450
rect 245120 443426 245148 452542
rect 245108 443420 245160 443426
rect 245108 443362 245160 443368
rect 242072 442332 242124 442338
rect 242072 442274 242124 442280
rect 242900 442332 242952 442338
rect 242900 442274 242952 442280
rect 242084 440298 242112 442274
rect 266372 440910 266400 697546
rect 282932 540258 282960 702406
rect 332520 700398 332548 703520
rect 332508 700392 332560 700398
rect 332508 700334 332560 700340
rect 348804 700330 348832 703520
rect 348792 700324 348844 700330
rect 348792 700266 348844 700272
rect 397472 699718 397500 703520
rect 397460 699712 397512 699718
rect 397460 699654 397512 699660
rect 403624 699712 403676 699718
rect 403624 699654 403676 699660
rect 403636 687206 403664 699654
rect 413664 698154 413692 703520
rect 462332 700369 462360 703520
rect 478524 700505 478552 703520
rect 478510 700496 478566 700505
rect 478510 700431 478566 700440
rect 462318 700360 462374 700369
rect 527192 700330 527220 703520
rect 543476 702434 543504 703520
rect 542372 702406 543504 702434
rect 462318 700295 462374 700304
rect 500224 700324 500276 700330
rect 500224 700266 500276 700272
rect 527180 700324 527232 700330
rect 527180 700266 527232 700272
rect 413652 698148 413704 698154
rect 413652 698090 413704 698096
rect 416044 698148 416096 698154
rect 416044 698090 416096 698096
rect 403624 687200 403676 687206
rect 403624 687142 403676 687148
rect 406384 687200 406436 687206
rect 406384 687142 406436 687148
rect 406396 647222 406424 687142
rect 416056 655518 416084 698090
rect 416044 655512 416096 655518
rect 416044 655454 416096 655460
rect 419448 655512 419500 655518
rect 419448 655454 419500 655460
rect 419460 651370 419488 655454
rect 419448 651364 419500 651370
rect 419448 651306 419500 651312
rect 424324 651364 424376 651370
rect 424324 651306 424376 651312
rect 406384 647216 406436 647222
rect 406384 647158 406436 647164
rect 409144 647216 409196 647222
rect 409144 647158 409196 647164
rect 409156 636886 409184 647158
rect 424336 638246 424364 651306
rect 424324 638240 424376 638246
rect 424324 638182 424376 638188
rect 432604 638240 432656 638246
rect 432604 638182 432656 638188
rect 409144 636880 409196 636886
rect 409144 636822 409196 636828
rect 414020 636880 414072 636886
rect 414020 636822 414072 636828
rect 414032 634098 414060 636822
rect 414020 634092 414072 634098
rect 414020 634034 414072 634040
rect 424140 634092 424192 634098
rect 424140 634034 424192 634040
rect 424152 628590 424180 634034
rect 424140 628584 424192 628590
rect 424140 628526 424192 628532
rect 432616 609278 432644 638182
rect 447784 628584 447836 628590
rect 447784 628526 447836 628532
rect 432604 609272 432656 609278
rect 432604 609214 432656 609220
rect 442264 609272 442316 609278
rect 442264 609214 442316 609220
rect 442276 579630 442304 609214
rect 447796 592006 447824 628526
rect 447784 592000 447836 592006
rect 447784 591942 447836 591948
rect 453304 592000 453356 592006
rect 453304 591942 453356 591948
rect 442264 579624 442316 579630
rect 442264 579566 442316 579572
rect 445668 579624 445720 579630
rect 445668 579566 445720 579572
rect 445680 574258 445708 579566
rect 445668 574252 445720 574258
rect 445668 574194 445720 574200
rect 447784 574252 447836 574258
rect 447784 574194 447836 574200
rect 447796 559774 447824 574194
rect 453316 562358 453344 591942
rect 453304 562352 453356 562358
rect 453304 562294 453356 562300
rect 456064 562352 456116 562358
rect 456064 562294 456116 562300
rect 447784 559768 447836 559774
rect 447784 559710 447836 559716
rect 451280 559768 451332 559774
rect 451280 559710 451332 559716
rect 451292 556850 451320 559710
rect 451280 556844 451332 556850
rect 451280 556786 451332 556792
rect 456076 554742 456104 562294
rect 461676 556844 461728 556850
rect 461676 556786 461728 556792
rect 461688 554742 461716 556786
rect 456064 554736 456116 554742
rect 456064 554678 456116 554684
rect 461584 554736 461636 554742
rect 461584 554678 461636 554684
rect 461676 554736 461728 554742
rect 461676 554678 461728 554684
rect 465724 554736 465776 554742
rect 465724 554678 465776 554684
rect 282920 540252 282972 540258
rect 282920 540194 282972 540200
rect 461596 538898 461624 554678
rect 461584 538892 461636 538898
rect 461584 538834 461636 538840
rect 465736 534750 465764 554678
rect 472624 538892 472676 538898
rect 472624 538834 472676 538840
rect 465724 534744 465776 534750
rect 465724 534686 465776 534692
rect 472636 529922 472664 538834
rect 475476 534744 475528 534750
rect 475476 534686 475528 534692
rect 472624 529916 472676 529922
rect 472624 529858 472676 529864
rect 475384 529916 475436 529922
rect 475384 529858 475436 529864
rect 475396 498817 475424 529858
rect 475488 526726 475516 534686
rect 475476 526720 475528 526726
rect 475476 526662 475528 526668
rect 479524 526720 479576 526726
rect 479524 526662 479576 526668
rect 479536 514078 479564 526662
rect 498844 524476 498896 524482
rect 498844 524418 498896 524424
rect 479524 514072 479576 514078
rect 479524 514014 479576 514020
rect 490564 514072 490616 514078
rect 490564 514014 490616 514020
rect 475382 498808 475438 498817
rect 475382 498743 475438 498752
rect 490576 488617 490604 514014
rect 490562 488608 490618 488617
rect 490562 488543 490618 488552
rect 266360 440904 266412 440910
rect 266360 440846 266412 440852
rect 240416 440292 240468 440298
rect 240416 440234 240468 440240
rect 242072 440292 242124 440298
rect 242072 440234 242124 440240
rect 240232 436620 240284 436626
rect 240232 436562 240284 436568
rect 240428 178906 240456 440234
rect 328196 180254 328348 180282
rect 335096 180254 335248 180282
rect 341996 180254 342148 180282
rect 366548 180260 366600 180266
rect 300124 180192 300176 180198
rect 241532 180118 241684 180146
rect 244752 180118 245088 180146
rect 248432 180118 248584 180146
rect 251192 180118 252080 180146
rect 255332 180118 255484 180146
rect 258092 180118 258980 180146
rect 262232 180118 262476 180146
rect 264992 180118 265880 180146
rect 269422 180118 269712 180146
rect 240416 178900 240468 178906
rect 240416 178842 240468 178848
rect 241532 177886 241560 180118
rect 241520 177880 241572 177886
rect 241520 177822 241572 177828
rect 244752 177342 244780 180118
rect 244740 177336 244792 177342
rect 244740 177278 244792 177284
rect 240048 177268 240100 177274
rect 240048 177210 240100 177216
rect 248432 60722 248460 180118
rect 248420 60716 248472 60722
rect 248420 60658 248472 60664
rect 251192 6798 251220 180118
rect 255332 100706 255360 180118
rect 255320 100700 255372 100706
rect 255320 100642 255372 100648
rect 258092 33114 258120 180118
rect 262232 139398 262260 180118
rect 262220 139392 262272 139398
rect 262220 139334 262272 139340
rect 264992 73166 265020 180118
rect 269684 177070 269712 180118
rect 271892 180118 272872 180146
rect 276322 180118 276704 180146
rect 269672 177064 269724 177070
rect 269672 177006 269724 177012
rect 271892 113150 271920 180118
rect 276676 177682 276704 180118
rect 278792 180118 279772 180146
rect 283314 180118 283696 180146
rect 286718 180118 286916 180146
rect 290214 180118 290504 180146
rect 293710 180118 293908 180146
rect 297114 180118 297496 180146
rect 300124 180134 300176 180140
rect 276664 177676 276716 177682
rect 276664 177618 276716 177624
rect 278792 153202 278820 180118
rect 283668 177614 283696 180118
rect 283656 177608 283708 177614
rect 283656 177550 283708 177556
rect 286888 176526 286916 180118
rect 290476 177410 290504 180118
rect 293880 177886 293908 180118
rect 295340 178832 295392 178838
rect 295340 178774 295392 178780
rect 293868 177880 293920 177886
rect 293868 177822 293920 177828
rect 290464 177404 290516 177410
rect 290464 177346 290516 177352
rect 286876 176520 286928 176526
rect 286876 176462 286928 176468
rect 295352 176254 295380 178774
rect 297468 177546 297496 180118
rect 300136 177886 300164 180134
rect 300610 180118 300808 180146
rect 304106 180118 304488 180146
rect 307510 180118 307708 180146
rect 311006 180118 311296 180146
rect 314502 180118 314608 180146
rect 317906 180118 318288 180146
rect 321402 180118 321508 180146
rect 324898 180118 325280 180146
rect 300124 177880 300176 177886
rect 300124 177822 300176 177828
rect 297456 177540 297508 177546
rect 297456 177482 297508 177488
rect 300780 176458 300808 180118
rect 304460 177478 304488 180118
rect 307680 178838 307708 180118
rect 307668 178832 307720 178838
rect 307668 178774 307720 178780
rect 311164 178764 311216 178770
rect 311164 178706 311216 178712
rect 304448 177472 304500 177478
rect 304448 177414 304500 177420
rect 300768 176452 300820 176458
rect 300768 176394 300820 176400
rect 295340 176248 295392 176254
rect 295340 176190 295392 176196
rect 311176 176186 311204 178706
rect 311268 176594 311296 180118
rect 311256 176588 311308 176594
rect 311256 176530 311308 176536
rect 314580 176390 314608 180118
rect 318260 178770 318288 180118
rect 318248 178764 318300 178770
rect 318248 178706 318300 178712
rect 321480 177206 321508 180118
rect 325252 179110 325280 180118
rect 325240 179104 325292 179110
rect 325240 179046 325292 179052
rect 328196 177886 328224 180254
rect 331798 180118 332088 180146
rect 328184 177880 328236 177886
rect 328184 177822 328236 177828
rect 332060 177313 332088 180118
rect 335096 179042 335124 180254
rect 338790 180118 339080 180146
rect 339052 179625 339080 180118
rect 339038 179616 339094 179625
rect 339038 179551 339094 179560
rect 335084 179036 335136 179042
rect 335084 178978 335136 178984
rect 341996 177818 342024 180254
rect 366548 180202 366600 180208
rect 367008 180260 367060 180266
rect 367008 180202 367060 180208
rect 345690 180118 346072 180146
rect 349186 180118 349568 180146
rect 352590 180118 352880 180146
rect 356086 180118 356376 180146
rect 359582 180118 359872 180146
rect 362986 180118 363368 180146
rect 346044 179722 346072 180118
rect 346032 179716 346084 179722
rect 346032 179658 346084 179664
rect 349540 178906 349568 180118
rect 348240 178900 348292 178906
rect 348240 178842 348292 178848
rect 349528 178900 349580 178906
rect 349528 178842 349580 178848
rect 348252 178022 348280 178842
rect 352852 178809 352880 180118
rect 352838 178800 352894 178809
rect 352838 178735 352894 178744
rect 348240 178016 348292 178022
rect 348240 177958 348292 177964
rect 356348 177857 356376 180118
rect 356334 177848 356390 177857
rect 341984 177812 342036 177818
rect 356334 177783 356390 177792
rect 341984 177754 342036 177760
rect 332046 177304 332102 177313
rect 332046 177239 332102 177248
rect 321468 177200 321520 177206
rect 321468 177142 321520 177148
rect 314568 176384 314620 176390
rect 314568 176326 314620 176332
rect 359844 176322 359872 180118
rect 363340 178498 363368 180118
rect 366100 180118 366436 180146
rect 363328 178492 363380 178498
rect 363328 178434 363380 178440
rect 359832 176316 359884 176322
rect 359832 176258 359884 176264
rect 366100 176186 366128 180118
rect 366560 177993 366588 180202
rect 366546 177984 366602 177993
rect 366546 177919 366602 177928
rect 367020 177313 367048 180202
rect 369978 180118 370360 180146
rect 370332 178673 370360 180118
rect 373000 180118 373336 180146
rect 376878 180118 377168 180146
rect 370318 178664 370374 178673
rect 370318 178599 370374 178608
rect 373000 178022 373028 180118
rect 372988 178016 373040 178022
rect 372988 177958 373040 177964
rect 377140 177342 377168 180118
rect 379992 180118 380328 180146
rect 383778 180118 383884 180146
rect 379992 177993 380020 180118
rect 380900 178696 380952 178702
rect 380900 178638 380952 178644
rect 380912 178022 380940 178638
rect 380992 178084 381044 178090
rect 380992 178026 381044 178032
rect 380900 178016 380952 178022
rect 379978 177984 380034 177993
rect 380900 177958 380952 177964
rect 379978 177919 380034 177928
rect 377128 177336 377180 177342
rect 367006 177304 367062 177313
rect 377128 177278 377180 177284
rect 367006 177239 367062 177248
rect 381004 177070 381032 178026
rect 380992 177064 381044 177070
rect 380992 177006 381044 177012
rect 383856 176254 383884 180118
rect 386892 180118 387228 180146
rect 390572 180118 390724 180146
rect 393792 180118 394128 180146
rect 397472 180118 397624 180146
rect 400784 180118 401120 180146
rect 404372 180118 404524 180146
rect 407684 180118 408020 180146
rect 411272 180118 411516 180146
rect 414676 180118 415012 180146
rect 418172 180118 418416 180146
rect 421576 180118 421912 180146
rect 425072 180118 425408 180146
rect 428476 180118 428812 180146
rect 432064 180118 432308 180146
rect 435272 180124 435324 180130
rect 386892 179858 386920 180118
rect 386880 179852 386932 179858
rect 386880 179794 386932 179800
rect 390572 177274 390600 180118
rect 393792 179586 393820 180118
rect 393780 179580 393832 179586
rect 393780 179522 393832 179528
rect 397472 178566 397500 180118
rect 398104 178696 398156 178702
rect 398104 178638 398156 178644
rect 397460 178560 397512 178566
rect 397460 178502 397512 178508
rect 390560 177268 390612 177274
rect 390560 177210 390612 177216
rect 398116 177206 398144 178638
rect 400784 177585 400812 180118
rect 404372 178634 404400 180118
rect 407684 179489 407712 180118
rect 407670 179480 407726 179489
rect 407670 179415 407726 179424
rect 411272 178945 411300 180118
rect 411258 178936 411314 178945
rect 411258 178871 411314 178880
rect 404360 178628 404412 178634
rect 404360 178570 404412 178576
rect 414676 178022 414704 180118
rect 418172 179081 418200 180118
rect 421576 179450 421604 180118
rect 421564 179444 421616 179450
rect 421564 179386 421616 179392
rect 425072 179217 425100 180118
rect 428476 179314 428504 180118
rect 432064 179790 432092 180118
rect 435272 180066 435324 180072
rect 435468 180118 435804 180146
rect 438872 180118 439208 180146
rect 442368 180118 442704 180146
rect 445864 180118 446200 180146
rect 449268 180118 449604 180146
rect 452764 180118 453100 180146
rect 455984 180118 456596 180146
rect 459664 180118 460000 180146
rect 463160 180118 463496 180146
rect 466656 180118 466992 180146
rect 470060 180118 470396 180146
rect 473556 180118 473892 180146
rect 477052 180118 477388 180146
rect 480548 180118 480792 180146
rect 483952 180118 484288 180146
rect 487172 180118 487784 180146
rect 489932 180118 491188 180146
rect 494072 180118 494684 180146
rect 498226 180118 498332 180146
rect 432052 179784 432104 179790
rect 432052 179726 432104 179732
rect 428464 179308 428516 179314
rect 428464 179250 428516 179256
rect 425058 179208 425114 179217
rect 425058 179143 425114 179152
rect 418158 179072 418214 179081
rect 418158 179007 418214 179016
rect 435284 178022 435312 180066
rect 414664 178016 414716 178022
rect 414664 177958 414716 177964
rect 435272 178016 435324 178022
rect 435272 177958 435324 177964
rect 435468 177721 435496 180118
rect 438872 179654 438900 180118
rect 438860 179648 438912 179654
rect 438860 179590 438912 179596
rect 435454 177712 435510 177721
rect 435454 177647 435510 177656
rect 400770 177576 400826 177585
rect 400770 177511 400826 177520
rect 442368 177449 442396 180118
rect 445864 179518 445892 180118
rect 445852 179512 445904 179518
rect 445852 179454 445904 179460
rect 449268 178022 449296 180118
rect 452764 179178 452792 180118
rect 452752 179172 452804 179178
rect 452752 179114 452804 179120
rect 449256 178016 449308 178022
rect 449256 177958 449308 177964
rect 455984 177750 456012 180118
rect 459664 179246 459692 180118
rect 459652 179240 459704 179246
rect 459652 179182 459704 179188
rect 463160 177954 463188 180118
rect 466656 179353 466684 180118
rect 466642 179344 466698 179353
rect 466642 179279 466698 179288
rect 463148 177948 463200 177954
rect 463148 177890 463200 177896
rect 455972 177744 456024 177750
rect 455972 177686 456024 177692
rect 456064 177744 456116 177750
rect 456064 177686 456116 177692
rect 442354 177440 442410 177449
rect 442354 177375 442410 177384
rect 398104 177200 398156 177206
rect 398104 177142 398156 177148
rect 383844 176248 383896 176254
rect 383844 176190 383896 176196
rect 311164 176180 311216 176186
rect 311164 176122 311216 176128
rect 366088 176180 366140 176186
rect 366088 176122 366140 176128
rect 278780 153196 278832 153202
rect 278780 153138 278832 153144
rect 456076 150414 456104 177686
rect 470060 177138 470088 180118
rect 473556 178974 473584 180118
rect 473544 178968 473596 178974
rect 473544 178910 473596 178916
rect 477052 177750 477080 180118
rect 477040 177744 477092 177750
rect 477040 177686 477092 177692
rect 470048 177132 470100 177138
rect 470048 177074 470100 177080
rect 480548 176662 480576 180118
rect 483952 179382 483980 180118
rect 483940 179376 483992 179382
rect 483940 179318 483992 179324
rect 483940 178968 483992 178974
rect 483940 178910 483992 178916
rect 485042 178936 485098 178945
rect 483952 177410 483980 178910
rect 485042 178871 485098 178880
rect 483940 177404 483992 177410
rect 483940 177346 483992 177352
rect 485056 177342 485084 178871
rect 485044 177336 485096 177342
rect 485044 177278 485096 177284
rect 480536 176656 480588 176662
rect 480536 176598 480588 176604
rect 456064 150408 456116 150414
rect 456064 150350 456116 150356
rect 487172 141438 487200 180118
rect 487160 141432 487212 141438
rect 487160 141374 487212 141380
rect 271880 113144 271932 113150
rect 271880 113086 271932 113092
rect 489932 85542 489960 180118
rect 492678 179480 492734 179489
rect 492678 179415 492734 179424
rect 492692 178226 492720 179415
rect 490932 178220 490984 178226
rect 490932 178162 490984 178168
rect 492680 178220 492732 178226
rect 492680 178162 492732 178168
rect 490944 176322 490972 178162
rect 493324 176724 493376 176730
rect 493324 176666 493376 176672
rect 490932 176316 490984 176322
rect 490932 176258 490984 176264
rect 489920 85536 489972 85542
rect 489920 85478 489972 85484
rect 264980 73160 265032 73166
rect 264980 73102 265032 73108
rect 258080 33108 258132 33114
rect 258080 33050 258132 33056
rect 493336 6866 493364 176666
rect 494072 45558 494100 180118
rect 498304 176730 498332 180118
rect 498856 178770 498884 524418
rect 499028 324352 499080 324358
rect 499028 324294 499080 324300
rect 499040 316034 499068 324294
rect 498948 316006 499068 316034
rect 498948 178838 498976 316006
rect 499028 271924 499080 271930
rect 499028 271866 499080 271872
rect 498936 178832 498988 178838
rect 498936 178774 498988 178780
rect 498844 178764 498896 178770
rect 498844 178706 498896 178712
rect 498292 176724 498344 176730
rect 498292 176666 498344 176672
rect 499040 176458 499068 271866
rect 499120 191888 499172 191894
rect 499120 191830 499172 191836
rect 499132 176526 499160 191830
rect 500236 178498 500264 700266
rect 501604 418192 501656 418198
rect 501604 418134 501656 418140
rect 500316 378208 500368 378214
rect 500316 378150 500368 378156
rect 500224 178492 500276 178498
rect 500224 178434 500276 178440
rect 499120 176520 499172 176526
rect 499120 176462 499172 176468
rect 499028 176452 499080 176458
rect 499028 176394 499080 176400
rect 500328 176390 500356 378150
rect 500408 258120 500460 258126
rect 500408 258062 500460 258068
rect 500420 177614 500448 258062
rect 500500 218068 500552 218074
rect 500500 218010 500552 218016
rect 500512 177682 500540 218010
rect 500500 177676 500552 177682
rect 500500 177618 500552 177624
rect 500408 177608 500460 177614
rect 500408 177550 500460 177556
rect 501616 177478 501644 418134
rect 501696 364404 501748 364410
rect 501696 364346 501748 364352
rect 501708 177546 501736 364346
rect 542372 179722 542400 702406
rect 580262 644056 580318 644065
rect 580262 643991 580318 644000
rect 580170 524512 580226 524521
rect 580170 524447 580172 524456
rect 580224 524447 580226 524456
rect 580172 524418 580224 524424
rect 580170 418296 580226 418305
rect 580170 418231 580226 418240
rect 580184 418198 580212 418231
rect 580172 418192 580224 418198
rect 580172 418134 580224 418140
rect 579802 378448 579858 378457
rect 579802 378383 579858 378392
rect 579816 378214 579844 378383
rect 579804 378208 579856 378214
rect 579804 378150 579856 378156
rect 580170 365120 580226 365129
rect 580170 365055 580226 365064
rect 580184 364410 580212 365055
rect 580172 364404 580224 364410
rect 580172 364346 580224 364352
rect 579986 325272 580042 325281
rect 579986 325207 580042 325216
rect 580000 324358 580028 325207
rect 579988 324352 580040 324358
rect 579988 324294 580040 324300
rect 580170 312080 580226 312089
rect 580170 312015 580226 312024
rect 579802 272232 579858 272241
rect 579802 272167 579858 272176
rect 579816 271930 579844 272167
rect 579804 271924 579856 271930
rect 579804 271866 579856 271872
rect 579986 258904 580042 258913
rect 579986 258839 580042 258848
rect 580000 258126 580028 258839
rect 579988 258120 580040 258126
rect 579988 258062 580040 258068
rect 580078 232384 580134 232393
rect 580078 232319 580134 232328
rect 579802 219056 579858 219065
rect 579802 218991 579858 219000
rect 579816 218074 579844 218991
rect 579804 218068 579856 218074
rect 579804 218010 579856 218016
rect 579986 192536 580042 192545
rect 579986 192471 580042 192480
rect 580000 191894 580028 192471
rect 579988 191888 580040 191894
rect 579988 191830 580040 191836
rect 580092 180198 580120 232319
rect 580080 180192 580132 180198
rect 580080 180134 580132 180140
rect 542360 179716 542412 179722
rect 542360 179658 542412 179664
rect 580184 179330 580212 312015
rect 580092 179302 580212 179330
rect 580092 178974 580120 179302
rect 580170 179208 580226 179217
rect 580170 179143 580226 179152
rect 580080 178968 580132 178974
rect 580080 178910 580132 178916
rect 580184 178090 580212 179143
rect 580276 178906 580304 643991
rect 580354 630864 580410 630873
rect 580354 630799 580410 630808
rect 580368 180266 580396 630799
rect 580446 591016 580502 591025
rect 580446 590951 580502 590960
rect 580356 180260 580408 180266
rect 580356 180202 580408 180208
rect 580264 178900 580316 178906
rect 580264 178842 580316 178848
rect 580172 178084 580224 178090
rect 580172 178026 580224 178032
rect 580460 177818 580488 590951
rect 580538 577688 580594 577697
rect 580538 577623 580594 577632
rect 580552 179110 580580 577623
rect 580630 537840 580686 537849
rect 580630 537775 580686 537784
rect 580540 179104 580592 179110
rect 580540 179046 580592 179052
rect 580644 179042 580672 537775
rect 580722 484664 580778 484673
rect 580722 484599 580778 484608
rect 580632 179036 580684 179042
rect 580632 178978 580684 178984
rect 580736 177886 580764 484599
rect 580814 471472 580870 471481
rect 580814 471407 580870 471416
rect 580828 185722 580856 471407
rect 580906 431624 580962 431633
rect 580906 431559 580962 431568
rect 580920 185842 580948 431559
rect 580908 185836 580960 185842
rect 580908 185778 580960 185784
rect 580828 185694 581040 185722
rect 580816 185632 580868 185638
rect 580816 185574 580868 185580
rect 580828 178702 580856 185574
rect 581012 185450 581040 185694
rect 580920 185422 581040 185450
rect 580816 178696 580868 178702
rect 580816 178638 580868 178644
rect 580724 177880 580776 177886
rect 580724 177822 580776 177828
rect 580448 177812 580500 177818
rect 580448 177754 580500 177760
rect 501696 177540 501748 177546
rect 501696 177482 501748 177488
rect 501604 177472 501656 177478
rect 501604 177414 501656 177420
rect 580920 176594 580948 185422
rect 580908 176588 580960 176594
rect 580908 176530 580960 176536
rect 500316 176384 500368 176390
rect 500316 176326 500368 176332
rect 580172 153196 580224 153202
rect 580172 153138 580224 153144
rect 580184 152697 580212 153138
rect 580170 152688 580226 152697
rect 580170 152623 580226 152632
rect 580172 139392 580224 139398
rect 580170 139360 580172 139369
rect 580224 139360 580226 139369
rect 580170 139295 580226 139304
rect 579804 113144 579856 113150
rect 579804 113086 579856 113092
rect 579816 112849 579844 113086
rect 579802 112840 579858 112849
rect 579802 112775 579858 112784
rect 580172 100700 580224 100706
rect 580172 100642 580224 100648
rect 580184 99521 580212 100642
rect 580170 99512 580226 99521
rect 580170 99447 580226 99456
rect 580172 73160 580224 73166
rect 580172 73102 580224 73108
rect 580184 73001 580212 73102
rect 580170 72992 580226 73001
rect 580170 72927 580226 72936
rect 580172 60716 580224 60722
rect 580172 60658 580224 60664
rect 580184 59673 580212 60658
rect 580170 59664 580226 59673
rect 580170 59599 580226 59608
rect 494060 45552 494112 45558
rect 494060 45494 494112 45500
rect 580170 33144 580226 33153
rect 580170 33079 580172 33088
rect 580224 33079 580226 33088
rect 580172 33050 580224 33056
rect 493324 6860 493376 6866
rect 493324 6802 493376 6808
rect 251180 6792 251232 6798
rect 251180 6734 251232 6740
rect 580172 6792 580224 6798
rect 580172 6734 580224 6740
rect 580184 6633 580212 6734
rect 580170 6624 580226 6633
rect 580170 6559 580226 6568
rect 47584 3460 47636 3466
rect 47584 3402 47636 3408
rect 1646 354 1758 480
rect 1412 326 1758 354
rect 1646 -960 1758 326
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 8114 700304 8170 700360
rect 3422 671200 3478 671256
rect 3422 658144 3478 658200
rect 3422 619112 3478 619168
rect 2870 501744 2926 501800
rect 2962 449520 3018 449576
rect 3330 397468 3332 397488
rect 3332 397468 3384 397488
rect 3384 397468 3386 397488
rect 3330 397432 3386 397468
rect 3146 306176 3202 306232
rect 3330 293120 3386 293176
rect 2778 254108 2834 254144
rect 2778 254088 2780 254108
rect 2780 254088 2832 254108
rect 2832 254088 2834 254108
rect 3146 241032 3202 241088
rect 2778 201864 2834 201920
rect 3514 606056 3570 606112
rect 3514 566888 3570 566944
rect 3606 553832 3662 553888
rect 3606 514800 3662 514856
rect 3698 462576 3754 462632
rect 3882 410488 3938 410544
rect 3790 358400 3846 358456
rect 3882 188808 3938 188864
rect 179418 465976 179474 466032
rect 91190 465160 91246 465216
rect 96158 465160 96214 465216
rect 98550 465160 98606 465216
rect 101678 465160 101734 465216
rect 103702 465160 103758 465216
rect 111062 465160 111118 465216
rect 113822 465160 113878 465216
rect 116214 465180 116270 465216
rect 116214 465160 116216 465180
rect 116216 465160 116268 465180
rect 116268 465160 116270 465180
rect 118606 465196 118608 465216
rect 118608 465196 118660 465216
rect 118660 465196 118662 465216
rect 118606 465160 118662 465196
rect 128726 465160 128782 465216
rect 136086 465160 136142 465216
rect 141054 465160 141110 465216
rect 143630 465160 143686 465216
rect 153382 465160 153438 465216
rect 156142 465160 156198 465216
rect 131118 463936 131174 463992
rect 168470 465160 168526 465216
rect 169758 465160 169814 465216
rect 83462 463664 83518 463720
rect 120998 463664 121054 463720
rect 123574 463664 123630 463720
rect 125966 463664 126022 463720
rect 133510 463664 133566 463720
rect 138478 463664 138534 463720
rect 146022 463664 146078 463720
rect 148506 463664 148562 463720
rect 151082 463664 151138 463720
rect 186870 465840 186926 465896
rect 188342 465704 188398 465760
rect 186870 461488 186926 461544
rect 7562 179424 7618 179480
rect 48042 416880 48098 416936
rect 47950 413752 48006 413808
rect 47582 388320 47638 388376
rect 47858 388048 47914 388104
rect 48134 415928 48190 415984
rect 49330 412800 49386 412856
rect 49238 409944 49294 410000
rect 48226 389952 48282 390008
rect 49422 411018 49478 411074
rect 49606 408162 49662 408218
rect 123482 379616 123538 379672
rect 130934 379616 130990 379672
rect 133510 379616 133566 379672
rect 145930 379616 145986 379672
rect 148506 379616 148562 379672
rect 155958 379616 156014 379672
rect 93950 379480 94006 379536
rect 96434 379480 96490 379536
rect 97630 379480 97686 379536
rect 98734 379480 98790 379536
rect 102230 379480 102286 379536
rect 125966 379480 126022 379536
rect 128542 379480 128598 379536
rect 150990 379208 151046 379264
rect 67546 377984 67602 378040
rect 73158 377984 73214 378040
rect 74354 377984 74410 378040
rect 78494 377984 78550 378040
rect 81162 377984 81218 378040
rect 92294 377984 92350 378040
rect 92846 377984 92902 378040
rect 95330 377984 95386 378040
rect 96526 377984 96582 378040
rect 99838 378020 99840 378040
rect 99840 378020 99892 378040
rect 99892 378020 99894 378040
rect 99838 377984 99894 378020
rect 101310 378004 101366 378040
rect 101310 377984 101312 378004
rect 101312 377984 101364 378004
rect 101364 377984 101366 378004
rect 66166 377032 66222 377088
rect 68926 377032 68982 377088
rect 70306 377032 70362 377088
rect 71686 377032 71742 377088
rect 73066 377032 73122 377088
rect 75826 377032 75882 377088
rect 77206 377032 77262 377088
rect 78310 377052 78366 377088
rect 78310 377032 78312 377052
rect 78312 377032 78364 377052
rect 78364 377032 78366 377052
rect 79966 377032 80022 377088
rect 81254 377032 81310 377088
rect 82726 377032 82782 377088
rect 84106 377032 84162 377088
rect 85486 377032 85542 377088
rect 86866 377032 86922 377088
rect 88154 377032 88210 377088
rect 89534 377032 89590 377088
rect 91006 377032 91062 377088
rect 91742 377052 91798 377088
rect 91742 377032 91744 377052
rect 91744 377032 91796 377052
rect 91796 377032 91798 377052
rect 81346 376896 81402 376952
rect 84014 376896 84070 376952
rect 86774 376896 86830 376952
rect 88246 376896 88302 376952
rect 89626 376896 89682 376952
rect 93766 377032 93822 377088
rect 103334 377984 103390 378040
rect 104806 377984 104862 378040
rect 105910 377984 105966 378040
rect 107566 377984 107622 378040
rect 110234 377984 110290 378040
rect 114466 377984 114522 378040
rect 120998 377984 121054 378040
rect 136086 377984 136142 378040
rect 139030 377984 139086 378040
rect 141606 377984 141662 378040
rect 143446 377984 143502 378040
rect 153382 377984 153438 378040
rect 104438 377868 104494 377904
rect 104438 377848 104440 377868
rect 104440 377848 104492 377868
rect 104492 377848 104494 377868
rect 99286 377032 99342 377088
rect 102046 377032 102102 377088
rect 106186 377032 106242 377088
rect 108946 377032 109002 377088
rect 111706 377032 111762 377088
rect 180706 377304 180762 377360
rect 117226 377032 117282 377088
rect 118606 377032 118662 377088
rect 173714 377032 173770 377088
rect 173806 376896 173862 376952
rect 49606 286320 49662 286376
rect 48134 236816 48190 236872
rect 47950 235864 48006 235920
rect 47858 233688 47914 233744
rect 47766 230968 47822 231024
rect 47674 229880 47730 229936
rect 47674 199008 47730 199064
rect 48042 232736 48098 232792
rect 47950 199824 48006 199880
rect 47858 199688 47914 199744
rect 49514 228162 49570 228218
rect 49330 209888 49386 209944
rect 48134 199552 48190 199608
rect 3422 149776 3478 149832
rect 3330 136720 3386 136776
rect 3146 84632 3202 84688
rect 3422 45500 3424 45520
rect 3424 45500 3476 45520
rect 3476 45500 3478 45520
rect 3422 45464 3478 45500
rect 3422 6432 3478 6488
rect 49422 208034 49478 208090
rect 136546 286220 136548 286240
rect 136548 286220 136600 286240
rect 136600 286220 136602 286240
rect 136546 286184 136602 286220
rect 139306 286184 139362 286240
rect 106186 285948 106188 285968
rect 106188 285948 106240 285968
rect 106240 285948 106242 285968
rect 106186 285912 106242 285948
rect 108946 285912 109002 285968
rect 144826 286184 144882 286240
rect 187698 465160 187754 465216
rect 187698 377304 187754 377360
rect 186962 376896 187018 376952
rect 189078 459176 189134 459232
rect 189078 399336 189134 399392
rect 189078 397704 189134 397760
rect 189262 396344 189318 396400
rect 189078 394848 189134 394904
rect 189262 393624 189318 393680
rect 180706 286320 180762 286376
rect 170678 286184 170734 286240
rect 83738 285676 83740 285696
rect 83740 285676 83792 285696
rect 83792 285676 83794 285696
rect 83738 285640 83794 285676
rect 86866 285640 86922 285696
rect 89626 285640 89682 285696
rect 92386 285660 92442 285696
rect 92386 285640 92388 285660
rect 92388 285640 92440 285660
rect 92440 285640 92442 285660
rect 93674 285640 93730 285696
rect 96526 285640 96582 285696
rect 104806 285640 104862 285696
rect 114466 285640 114522 285696
rect 118606 285640 118662 285696
rect 124126 285640 124182 285696
rect 126886 285640 126942 285696
rect 133786 285640 133842 285696
rect 141882 285640 141938 285696
rect 151726 285640 151782 285696
rect 154486 285640 154542 285696
rect 157246 285640 157302 285696
rect 169666 285640 169722 285696
rect 128726 285132 128728 285152
rect 128728 285132 128780 285152
rect 128780 285132 128782 285152
rect 128726 285096 128782 285132
rect 131118 285096 131174 285152
rect 111062 284996 111064 285016
rect 111064 284996 111116 285016
rect 111116 284996 111118 285016
rect 111062 284960 111118 284996
rect 116214 284960 116270 285016
rect 98550 284824 98606 284880
rect 148598 284860 148600 284880
rect 148600 284860 148652 284880
rect 148652 284860 148654 284880
rect 148598 284824 148654 284860
rect 101310 284688 101366 284744
rect 146022 284724 146024 284744
rect 146024 284724 146076 284744
rect 146076 284724 146078 284744
rect 146022 284688 146078 284724
rect 180706 284008 180762 284064
rect 49606 208306 49662 208362
rect 71870 199416 71926 199472
rect 77758 199416 77814 199472
rect 81346 199416 81402 199472
rect 82542 199416 82598 199472
rect 83462 199416 83518 199472
rect 86222 199416 86278 199472
rect 103702 199436 103758 199472
rect 103702 199416 103704 199436
rect 103704 199416 103756 199436
rect 103756 199416 103758 199436
rect 70582 198600 70638 198656
rect 76654 198600 76710 198656
rect 78862 198600 78918 198656
rect 80150 198600 80206 198656
rect 84566 198636 84568 198656
rect 84568 198636 84620 198656
rect 84620 198636 84622 198656
rect 84566 198600 84622 198636
rect 88246 198620 88302 198656
rect 88246 198600 88248 198620
rect 88248 198600 88300 198620
rect 88300 198600 88302 198620
rect 67546 198192 67602 198248
rect 66166 197376 66222 197432
rect 74354 198192 74410 198248
rect 88614 198600 88670 198656
rect 91190 198600 91246 198656
rect 93582 198600 93638 198656
rect 93950 198600 94006 198656
rect 95974 198600 96030 198656
rect 98366 198600 98422 198656
rect 99838 198600 99894 198656
rect 100942 198600 100998 198656
rect 102230 198600 102286 198656
rect 85854 198464 85910 198520
rect 87418 198464 87474 198520
rect 90914 198464 90970 198520
rect 68926 197376 68982 197432
rect 69846 197376 69902 197432
rect 75734 198056 75790 198112
rect 74446 197376 74502 197432
rect 83738 197920 83794 197976
rect 78586 197376 78642 197432
rect 81070 197376 81126 197432
rect 89534 198328 89590 198384
rect 92846 198328 92902 198384
rect 92294 198192 92350 198248
rect 128358 199280 128414 199336
rect 106094 198600 106150 198656
rect 107014 198600 107070 198656
rect 108486 198600 108542 198656
rect 113638 198600 113694 198656
rect 120998 198600 121054 198656
rect 123574 198600 123630 198656
rect 105910 197920 105966 197976
rect 111062 197920 111118 197976
rect 116214 197784 116270 197840
rect 118422 197784 118478 197840
rect 128542 198600 128598 198656
rect 130934 198600 130990 198656
rect 136086 198600 136142 198656
rect 150990 199416 151046 199472
rect 138754 198600 138810 198656
rect 143446 198600 143502 198656
rect 146022 198600 146078 198656
rect 148598 198600 148654 198656
rect 153382 198600 153438 198656
rect 173438 198600 173494 198656
rect 126150 197648 126206 197704
rect 133510 197648 133566 197704
rect 138754 196832 138810 196888
rect 143446 196696 143502 196752
rect 155958 197784 156014 197840
rect 173254 197784 173310 197840
rect 187146 198464 187202 198520
rect 187606 205672 187662 205728
rect 187330 198328 187386 198384
rect 189078 219272 189134 219328
rect 189078 216280 189134 216336
rect 189998 279112 190054 279168
rect 189906 217640 189962 217696
rect 190090 214784 190146 214840
rect 190274 213560 190330 213616
rect 191194 379344 191250 379400
rect 195242 465568 195298 465624
rect 232502 285776 232558 285832
rect 237470 438096 237526 438152
rect 237378 437552 237434 437608
rect 237470 433608 237526 433664
rect 237378 433372 237380 433392
rect 237380 433372 237432 433392
rect 237432 433372 237434 433392
rect 237378 433336 237434 433372
rect 237378 431296 237434 431352
rect 237378 429256 237434 429312
rect 237378 428440 237434 428496
rect 237378 426264 237434 426320
rect 237378 425176 237434 425232
rect 237378 423952 237434 424008
rect 237378 422048 237434 422104
rect 237378 420980 237434 421016
rect 237378 420960 237380 420980
rect 237380 420960 237432 420980
rect 237432 420960 237434 420980
rect 237378 419600 237434 419656
rect 237470 416064 237526 416120
rect 237378 415520 237434 415576
rect 237378 413752 237434 413808
rect 237378 411712 237434 411768
rect 237378 407360 237434 407416
rect 237378 405048 237434 405104
rect 237378 403280 237434 403336
rect 237378 400016 237434 400072
rect 237378 398928 237434 398984
rect 237378 395972 237380 395992
rect 237380 395972 237432 395992
rect 237432 395972 237434 395992
rect 237378 395936 237434 395972
rect 237378 394732 237434 394768
rect 237378 394712 237380 394732
rect 237380 394712 237432 394732
rect 237432 394712 237434 394732
rect 237378 391892 237380 391912
rect 237380 391892 237432 391912
rect 237432 391892 237434 391912
rect 237378 391856 237434 391892
rect 237470 389680 237526 389736
rect 237378 389272 237434 389328
rect 237378 387368 237434 387424
rect 237378 385328 237434 385384
rect 237470 385056 237526 385112
rect 237378 383016 237434 383072
rect 237378 380976 237434 381032
rect 237378 380024 237434 380080
rect 237378 377304 237434 377360
rect 237378 376660 237380 376680
rect 237380 376660 237432 376680
rect 237432 376660 237434 376680
rect 237378 376624 237434 376660
rect 237378 373360 237434 373416
rect 237378 372272 237434 372328
rect 237378 368364 237380 368384
rect 237380 368364 237432 368384
rect 237432 368364 237434 368384
rect 237378 368328 237434 368364
rect 237470 368056 237526 368112
rect 238574 440136 238630 440192
rect 238482 435784 238538 435840
rect 238390 418104 238446 418160
rect 238390 411304 238446 411360
rect 238298 409400 238354 409456
rect 238298 406408 238354 406464
rect 238482 402056 238538 402112
rect 238574 397568 238630 397624
rect 238666 393352 238722 393408
rect 238206 373904 238262 373960
rect 238114 369688 238170 369744
rect 238022 365472 238078 365528
rect 237378 364112 237434 364168
rect 237470 363704 237526 363760
rect 237378 361120 237434 361176
rect 237378 359896 237434 359952
rect 237378 358708 237380 358728
rect 237380 358708 237432 358728
rect 237432 358708 237434 358728
rect 237378 358672 237434 358708
rect 237378 355816 237434 355872
rect 237378 354628 237380 354648
rect 237380 354628 237432 354648
rect 237432 354628 237434 354648
rect 237378 354592 237434 354628
rect 237378 351464 237434 351520
rect 237378 350240 237434 350296
rect 237378 347520 237434 347576
rect 237470 346976 237526 347032
rect 237378 346160 237434 346216
rect 237378 343440 237434 343496
rect 237378 342116 237380 342136
rect 237380 342116 237432 342136
rect 237432 342116 237434 342136
rect 237378 342080 237434 342116
rect 237470 341808 237526 341864
rect 237378 339088 237434 339144
rect 237378 337864 237434 337920
rect 237470 337320 237526 337376
rect 237378 336504 237434 336560
rect 237378 335144 237434 335200
rect 237470 334736 237526 334792
rect 237378 333784 237434 333840
rect 237378 332424 237434 332480
rect 237470 332152 237526 332208
rect 237378 330928 237434 330984
rect 237378 329432 237434 329488
rect 237378 328208 237434 328264
rect 237470 327664 237526 327720
rect 237378 326848 237434 326904
rect 237470 325524 237472 325544
rect 237472 325524 237524 325544
rect 237524 325524 237526 325544
rect 237470 325488 237526 325524
rect 237378 325080 237434 325136
rect 237378 324128 237434 324184
rect 237378 322768 237434 322824
rect 237378 321408 237434 321464
rect 237378 320068 237434 320104
rect 237378 320048 237380 320068
rect 237380 320048 237432 320068
rect 237432 320048 237434 320068
rect 237470 319776 237526 319832
rect 237378 318552 237434 318608
rect 238298 322360 238354 322416
rect 238022 318008 238078 318064
rect 237378 317192 237434 317248
rect 237378 315424 237434 315480
rect 237378 314472 237434 314528
rect 237378 313148 237380 313168
rect 237380 313148 237432 313168
rect 237432 313148 237434 313168
rect 237378 313112 237434 313148
rect 237470 312704 237526 312760
rect 237378 311788 237380 311808
rect 237380 311788 237432 311808
rect 237432 311788 237434 311808
rect 237378 311752 237434 311788
rect 237378 310412 237434 310448
rect 237378 310392 237380 310412
rect 237380 310392 237432 310412
rect 237432 310392 237434 310412
rect 237470 310120 237526 310176
rect 237378 308896 237434 308952
rect 237470 308352 237526 308408
rect 237378 307536 237434 307592
rect 237378 306176 237434 306232
rect 237470 305768 237526 305824
rect 237378 304816 237434 304872
rect 237378 303456 237434 303512
rect 237470 303048 237526 303104
rect 237378 302132 237380 302152
rect 237380 302132 237432 302152
rect 237432 302132 237434 302152
rect 237378 302096 237434 302132
rect 237378 300772 237380 300792
rect 237380 300772 237432 300792
rect 237432 300772 237434 300792
rect 237378 300736 237434 300772
rect 237470 300464 237526 300520
rect 237378 299240 237434 299296
rect 237470 298696 237526 298752
rect 237378 297880 237434 297936
rect 237378 296520 237434 296576
rect 237470 296112 237526 296168
rect 237378 295160 237434 295216
rect 237378 293800 237434 293856
rect 237378 292712 237434 292768
rect 234986 199688 235042 199744
rect 235170 199552 235226 199608
rect 235446 197104 235502 197160
rect 233974 179152 234030 179208
rect 237378 291352 237434 291408
rect 237378 289992 237434 290048
rect 237470 288632 237526 288688
rect 237378 288496 237434 288552
rect 237378 287136 237434 287192
rect 237378 286048 237434 286104
rect 237470 285796 237526 285832
rect 237470 285776 237472 285796
rect 237472 285776 237524 285796
rect 237524 285776 237526 285796
rect 237378 284860 237380 284880
rect 237380 284860 237432 284880
rect 237432 284860 237434 284880
rect 237378 284824 237434 284860
rect 237378 283464 237434 283520
rect 237470 282940 237526 282976
rect 237470 282920 237472 282940
rect 237472 282920 237524 282940
rect 237524 282920 237526 282940
rect 237378 282820 237380 282840
rect 237380 282820 237432 282840
rect 237432 282820 237434 282840
rect 237378 282784 237434 282820
rect 237378 280744 237434 280800
rect 237470 280336 237526 280392
rect 237378 279792 237434 279848
rect 237378 277208 237434 277264
rect 237470 275032 237526 275088
rect 237378 274488 237434 274544
rect 237378 271804 237380 271824
rect 237380 271804 237432 271824
rect 237432 271804 237434 271824
rect 237378 271768 237434 271804
rect 237838 269728 237894 269784
rect 237378 267824 237434 267880
rect 237378 262384 237434 262440
rect 237378 261976 237434 262032
rect 237470 261840 237526 261896
rect 237378 259664 237434 259720
rect 237470 259528 237526 259584
rect 237378 259120 237434 259176
rect 237378 257080 237434 257136
rect 237470 256828 237526 256864
rect 237470 256808 237472 256828
rect 237472 256808 237524 256828
rect 237524 256808 237526 256828
rect 237470 254496 237526 254552
rect 237378 254088 237434 254144
rect 237378 251776 237434 251832
rect 237378 249872 237434 249928
rect 237378 248512 237434 248568
rect 237378 247052 237380 247072
rect 237380 247052 237432 247072
rect 237432 247052 237434 247072
rect 237378 247016 237434 247052
rect 237378 244432 237434 244488
rect 237378 242836 237380 242856
rect 237380 242836 237432 242856
rect 237432 242836 237434 242856
rect 237378 242800 237434 242836
rect 237378 241576 237434 241632
rect 237378 240352 237434 240408
rect 237378 238584 237434 238640
rect 237378 236020 237434 236056
rect 237378 236000 237380 236020
rect 237380 236000 237432 236020
rect 237432 236000 237434 236020
rect 237378 234232 237434 234288
rect 237378 232464 237434 232520
rect 237378 230152 237434 230208
rect 237470 228112 237526 228168
rect 237378 227740 237380 227760
rect 237380 227740 237432 227760
rect 237432 227740 237434 227760
rect 237378 227704 237434 227740
rect 238114 253816 238170 253872
rect 238114 251368 238170 251424
rect 238022 225800 238078 225856
rect 237378 223644 237434 223680
rect 237378 223624 237380 223644
rect 237380 223624 237432 223644
rect 237432 223624 237434 223644
rect 237470 222808 237526 222864
rect 237378 222284 237434 222320
rect 237378 222264 237380 222284
rect 237380 222264 237432 222284
rect 237432 222264 237434 222284
rect 237470 221584 237526 221640
rect 237378 221448 237434 221504
rect 237378 219544 237434 219600
rect 237470 218456 237526 218512
rect 237378 218084 237380 218104
rect 237380 218084 237432 218104
rect 237432 218084 237434 218104
rect 237378 218048 237434 218084
rect 237378 216416 237434 216472
rect 238022 215328 238078 215384
rect 237378 213424 237434 213480
rect 237470 212744 237526 212800
rect 237378 212336 237434 212392
rect 237470 209888 237526 209944
rect 237378 209616 237434 209672
rect 237378 208412 237434 208448
rect 237378 208392 237380 208412
rect 237380 208392 237432 208412
rect 237432 208392 237434 208412
rect 237470 208292 237472 208312
rect 237472 208292 237524 208312
rect 237524 208292 237526 208312
rect 237470 208256 237526 208292
rect 237930 206080 237986 206136
rect 237470 205808 237526 205864
rect 237378 205572 237380 205592
rect 237380 205572 237432 205592
rect 237432 205572 237434 205592
rect 237378 205536 237434 205572
rect 237378 203496 237434 203552
rect 237470 202952 237526 203008
rect 237378 202544 237434 202600
rect 237378 201492 237380 201512
rect 237380 201492 237432 201512
rect 237432 201492 237434 201512
rect 237378 201456 237434 201492
rect 237470 200096 237526 200152
rect 237378 199960 237434 200016
rect 237378 197956 237380 197976
rect 237380 197956 237432 197976
rect 237432 197956 237434 197976
rect 237378 197920 237434 197956
rect 237378 197276 237380 197296
rect 237380 197276 237432 197296
rect 237432 197276 237434 197296
rect 237378 197240 237434 197276
rect 238298 270680 238354 270736
rect 238206 248240 238262 248296
rect 238206 245656 238262 245712
rect 238482 267144 238538 267200
rect 238482 264968 238538 265024
rect 238390 245520 238446 245576
rect 238390 243072 238446 243128
rect 238298 213968 238354 214024
rect 238666 264016 238722 264072
rect 238574 250824 238630 250880
rect 238574 237360 238630 237416
rect 238482 211112 238538 211168
rect 238666 232056 238722 232112
rect 237470 196036 237526 196072
rect 237470 196016 237472 196036
rect 237472 196016 237524 196036
rect 237524 196016 237526 196036
rect 237378 195916 237380 195936
rect 237380 195916 237432 195936
rect 237432 195916 237434 195936
rect 237378 195880 237434 195916
rect 237378 194420 237380 194440
rect 237380 194420 237432 194440
rect 237432 194420 237434 194440
rect 237378 194384 237434 194420
rect 237470 194112 237526 194168
rect 237378 192888 237434 192944
rect 237470 191700 237472 191720
rect 237472 191700 237524 191720
rect 237524 191700 237526 191720
rect 237470 191664 237526 191700
rect 237378 191528 237434 191584
rect 237378 190304 237434 190360
rect 237470 189760 237526 189816
rect 237378 188980 237380 189000
rect 237380 188980 237432 189000
rect 237432 188980 237434 189000
rect 237378 188944 237434 188980
rect 237378 187620 237380 187640
rect 237380 187620 237432 187640
rect 237432 187620 237434 187640
rect 237378 187584 237434 187620
rect 237378 186260 237380 186280
rect 237380 186260 237432 186280
rect 237432 186260 237434 186280
rect 237378 186224 237434 186260
rect 237378 184884 237434 184920
rect 237378 184864 237380 184884
rect 237380 184864 237432 184884
rect 237432 184864 237434 184884
rect 237470 184456 237526 184512
rect 237378 183232 237434 183288
rect 237378 182008 237434 182064
rect 237470 181872 237526 181928
rect 237562 180648 237618 180704
rect 239494 178880 239550 178936
rect 238758 177656 238814 177712
rect 237378 177520 237434 177576
rect 191194 177384 191250 177440
rect 478510 700440 478566 700496
rect 462318 700304 462374 700360
rect 475382 498752 475438 498808
rect 490562 488552 490618 488608
rect 339038 179560 339094 179616
rect 352838 178744 352894 178800
rect 356334 177792 356390 177848
rect 332046 177248 332102 177304
rect 366546 177928 366602 177984
rect 370318 178608 370374 178664
rect 379978 177928 380034 177984
rect 367006 177248 367062 177304
rect 407670 179424 407726 179480
rect 411258 178880 411314 178936
rect 425058 179152 425114 179208
rect 418158 179016 418214 179072
rect 435454 177656 435510 177712
rect 400770 177520 400826 177576
rect 466642 179288 466698 179344
rect 442354 177384 442410 177440
rect 485042 178880 485098 178936
rect 492678 179424 492734 179480
rect 580262 644000 580318 644056
rect 580170 524476 580226 524512
rect 580170 524456 580172 524476
rect 580172 524456 580224 524476
rect 580224 524456 580226 524476
rect 580170 418240 580226 418296
rect 579802 378392 579858 378448
rect 580170 365064 580226 365120
rect 579986 325216 580042 325272
rect 580170 312024 580226 312080
rect 579802 272176 579858 272232
rect 579986 258848 580042 258904
rect 580078 232328 580134 232384
rect 579802 219000 579858 219056
rect 579986 192480 580042 192536
rect 580170 179152 580226 179208
rect 580354 630808 580410 630864
rect 580446 590960 580502 591016
rect 580538 577632 580594 577688
rect 580630 537784 580686 537840
rect 580722 484608 580778 484664
rect 580814 471416 580870 471472
rect 580906 431568 580962 431624
rect 580170 152632 580226 152688
rect 580170 139340 580172 139360
rect 580172 139340 580224 139360
rect 580224 139340 580226 139360
rect 580170 139304 580226 139340
rect 579802 112784 579858 112840
rect 580170 99456 580226 99512
rect 580170 72936 580226 72992
rect 580170 59608 580226 59664
rect 580170 33108 580226 33144
rect 580170 33088 580172 33108
rect 580172 33088 580224 33108
rect 580224 33088 580226 33108
rect 580170 6568 580226 6624
<< metal3 >>
rect 478505 700498 478571 700501
rect 491334 700498 491340 700500
rect 478505 700496 491340 700498
rect 478505 700440 478510 700496
rect 478566 700440 491340 700496
rect 478505 700438 491340 700440
rect 478505 700435 478571 700438
rect 491334 700436 491340 700438
rect 491404 700436 491410 700500
rect 8109 700362 8175 700365
rect 239254 700362 239260 700364
rect 8109 700360 239260 700362
rect 8109 700304 8114 700360
rect 8170 700304 239260 700360
rect 8109 700302 239260 700304
rect 8109 700299 8175 700302
rect 239254 700300 239260 700302
rect 239324 700300 239330 700364
rect 462313 700362 462379 700365
rect 492806 700362 492812 700364
rect 462313 700360 492812 700362
rect 462313 700304 462318 700360
rect 462374 700304 492812 700360
rect 462313 700302 492812 700304
rect 462313 700299 462379 700302
rect 492806 700300 492812 700302
rect 492876 700300 492882 700364
rect -960 697220 480 697460
rect 580206 697172 580212 697236
rect 580276 697234 580282 697236
rect 583520 697234 584960 697324
rect 580276 697174 584960 697234
rect 580276 697172 580282 697174
rect 583520 697084 584960 697174
rect -960 684164 480 684404
rect 580390 683844 580396 683908
rect 580460 683906 580466 683908
rect 583520 683906 584960 683996
rect 580460 683846 584960 683906
rect 580460 683844 580466 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3417 671258 3483 671261
rect -960 671256 3483 671258
rect -960 671200 3422 671256
rect 3478 671200 3483 671256
rect -960 671198 3483 671200
rect -960 671108 480 671198
rect 3417 671195 3483 671198
rect 583520 670564 584960 670804
rect -960 658202 480 658292
rect 3417 658202 3483 658205
rect -960 658200 3483 658202
rect -960 658144 3422 658200
rect 3478 658144 3483 658200
rect -960 658142 3483 658144
rect -960 658052 480 658142
rect 3417 658139 3483 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 580257 644058 580323 644061
rect 583520 644058 584960 644148
rect 580257 644056 584960 644058
rect 580257 644000 580262 644056
rect 580318 644000 584960 644056
rect 580257 643998 584960 644000
rect 580257 643995 580323 643998
rect 583520 643908 584960 643998
rect -960 631940 480 632180
rect 580349 630866 580415 630869
rect 583520 630866 584960 630956
rect 580349 630864 584960 630866
rect 580349 630808 580354 630864
rect 580410 630808 584960 630864
rect 580349 630806 584960 630808
rect 580349 630803 580415 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3417 619170 3483 619173
rect -960 619168 3483 619170
rect -960 619112 3422 619168
rect 3478 619112 3483 619168
rect -960 619110 3483 619112
rect -960 619020 480 619110
rect 3417 619107 3483 619110
rect 583520 617388 584960 617628
rect -960 606114 480 606204
rect 3509 606114 3575 606117
rect -960 606112 3575 606114
rect -960 606056 3514 606112
rect 3570 606056 3575 606112
rect -960 606054 3575 606056
rect -960 605964 480 606054
rect 3509 606051 3575 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 580441 591018 580507 591021
rect 583520 591018 584960 591108
rect 580441 591016 584960 591018
rect 580441 590960 580446 591016
rect 580502 590960 584960 591016
rect 580441 590958 584960 590960
rect 580441 590955 580507 590958
rect 583520 590868 584960 590958
rect -960 579852 480 580092
rect 580533 577690 580599 577693
rect 583520 577690 584960 577780
rect 580533 577688 584960 577690
rect 580533 577632 580538 577688
rect 580594 577632 584960 577688
rect 580533 577630 584960 577632
rect 580533 577627 580599 577630
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 3509 566946 3575 566949
rect -960 566944 3575 566946
rect -960 566888 3514 566944
rect 3570 566888 3575 566944
rect -960 566886 3575 566888
rect -960 566796 480 566886
rect 3509 566883 3575 566886
rect 583520 564212 584960 564452
rect -960 553890 480 553980
rect 3601 553890 3667 553893
rect -960 553888 3667 553890
rect -960 553832 3606 553888
rect 3662 553832 3667 553888
rect -960 553830 3667 553832
rect -960 553740 480 553830
rect 3601 553827 3667 553830
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 580625 537842 580691 537845
rect 583520 537842 584960 537932
rect 580625 537840 584960 537842
rect 580625 537784 580630 537840
rect 580686 537784 584960 537840
rect 580625 537782 584960 537784
rect 580625 537779 580691 537782
rect 583520 537692 584960 537782
rect -960 527764 480 528004
rect 580165 524514 580231 524517
rect 583520 524514 584960 524604
rect 580165 524512 584960 524514
rect 580165 524456 580170 524512
rect 580226 524456 584960 524512
rect 580165 524454 584960 524456
rect 580165 524451 580231 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 3601 514858 3667 514861
rect -960 514856 3667 514858
rect -960 514800 3606 514856
rect 3662 514800 3667 514856
rect -960 514798 3667 514800
rect -960 514708 480 514798
rect 3601 514795 3667 514798
rect 583520 511172 584960 511412
rect -960 501802 480 501892
rect 2865 501802 2931 501805
rect -960 501800 2931 501802
rect -960 501744 2870 501800
rect 2926 501744 2931 501800
rect -960 501742 2931 501744
rect -960 501652 480 501742
rect 2865 501739 2931 501742
rect 475377 498810 475443 498813
rect 490414 498810 490420 498812
rect 475377 498808 490420 498810
rect 475377 498752 475382 498808
rect 475438 498752 490420 498808
rect 475377 498750 490420 498752
rect 475377 498747 475443 498750
rect 490414 498748 490420 498750
rect 490484 498748 490490 498812
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 490557 488610 490623 488613
rect 494094 488610 494100 488612
rect 490557 488608 494100 488610
rect 490557 488552 490562 488608
rect 490618 488552 494100 488608
rect 490557 488550 494100 488552
rect 490557 488547 490623 488550
rect 494094 488548 494100 488550
rect 494164 488548 494170 488612
rect 580717 484666 580783 484669
rect 583520 484666 584960 484756
rect 580717 484664 584960 484666
rect 580717 484608 580722 484664
rect 580778 484608 584960 484664
rect 580717 484606 584960 484608
rect 580717 484603 580783 484606
rect 583520 484516 584960 484606
rect -960 475540 480 475780
rect 580809 471474 580875 471477
rect 583520 471474 584960 471564
rect 580809 471472 584960 471474
rect 580809 471416 580814 471472
rect 580870 471416 584960 471472
rect 580809 471414 584960 471416
rect 580809 471411 580875 471414
rect 583520 471324 584960 471414
rect 86166 466108 86172 466172
rect 86236 466170 86242 466172
rect 237966 466170 237972 466172
rect 86236 466110 237972 466170
rect 86236 466108 86242 466110
rect 237966 466108 237972 466110
rect 238036 466108 238042 466172
rect 88558 465972 88564 466036
rect 88628 466034 88634 466036
rect 179413 466034 179479 466037
rect 88628 466032 179479 466034
rect 88628 465976 179418 466032
rect 179474 465976 179479 466032
rect 88628 465974 179479 465976
rect 88628 465972 88634 465974
rect 179413 465971 179479 465974
rect 93526 465836 93532 465900
rect 93596 465898 93602 465900
rect 186865 465898 186931 465901
rect 93596 465896 186931 465898
rect 93596 465840 186870 465896
rect 186926 465840 186931 465896
rect 93596 465838 186931 465840
rect 93596 465836 93602 465838
rect 186865 465835 186931 465838
rect 81014 465700 81020 465764
rect 81084 465762 81090 465764
rect 188337 465762 188403 465765
rect 81084 465760 188403 465762
rect 81084 465704 188342 465760
rect 188398 465704 188403 465760
rect 81084 465702 188403 465704
rect 81084 465700 81090 465702
rect 188337 465699 188403 465702
rect 78806 465564 78812 465628
rect 78876 465626 78882 465628
rect 195237 465626 195303 465629
rect 78876 465624 195303 465626
rect 78876 465568 195242 465624
rect 195298 465568 195303 465624
rect 78876 465566 195303 465568
rect 78876 465564 78882 465566
rect 195237 465563 195303 465566
rect 108430 465428 108436 465492
rect 108500 465490 108506 465492
rect 238518 465490 238524 465492
rect 108500 465430 238524 465490
rect 108500 465428 108506 465430
rect 238518 465428 238524 465430
rect 238588 465428 238594 465492
rect 106222 465292 106228 465356
rect 106292 465354 106298 465356
rect 238334 465354 238340 465356
rect 106292 465294 238340 465354
rect 106292 465292 106298 465294
rect 238334 465292 238340 465294
rect 238404 465292 238410 465356
rect 91185 465220 91251 465221
rect 96153 465220 96219 465221
rect 98545 465220 98611 465221
rect 91134 465218 91140 465220
rect 91094 465158 91140 465218
rect 91204 465216 91251 465220
rect 96102 465218 96108 465220
rect 91246 465160 91251 465216
rect 91134 465156 91140 465158
rect 91204 465156 91251 465160
rect 96062 465158 96108 465218
rect 96172 465216 96219 465220
rect 98494 465218 98500 465220
rect 96214 465160 96219 465216
rect 96102 465156 96108 465158
rect 96172 465156 96219 465160
rect 98454 465158 98500 465218
rect 98564 465216 98611 465220
rect 98606 465160 98611 465216
rect 98494 465156 98500 465158
rect 98564 465156 98611 465160
rect 101254 465156 101260 465220
rect 101324 465218 101330 465220
rect 101673 465218 101739 465221
rect 103697 465220 103763 465221
rect 111057 465220 111123 465221
rect 113817 465220 113883 465221
rect 116209 465220 116275 465221
rect 118601 465220 118667 465221
rect 128721 465220 128787 465221
rect 136081 465220 136147 465221
rect 141049 465220 141115 465221
rect 143625 465220 143691 465221
rect 153377 465220 153443 465221
rect 156137 465220 156203 465221
rect 168465 465220 168531 465221
rect 169753 465220 169819 465221
rect 103646 465218 103652 465220
rect 101324 465216 101739 465218
rect 101324 465160 101678 465216
rect 101734 465160 101739 465216
rect 101324 465158 101739 465160
rect 103606 465158 103652 465218
rect 103716 465216 103763 465220
rect 111006 465218 111012 465220
rect 103758 465160 103763 465216
rect 101324 465156 101330 465158
rect 91185 465155 91251 465156
rect 96153 465155 96219 465156
rect 98545 465155 98611 465156
rect 101673 465155 101739 465158
rect 103646 465156 103652 465158
rect 103716 465156 103763 465160
rect 110966 465158 111012 465218
rect 111076 465216 111123 465220
rect 113766 465218 113772 465220
rect 111118 465160 111123 465216
rect 111006 465156 111012 465158
rect 111076 465156 111123 465160
rect 113726 465158 113772 465218
rect 113836 465216 113883 465220
rect 116158 465218 116164 465220
rect 113878 465160 113883 465216
rect 113766 465156 113772 465158
rect 113836 465156 113883 465160
rect 116118 465158 116164 465218
rect 116228 465216 116275 465220
rect 118550 465218 118556 465220
rect 116270 465160 116275 465216
rect 116158 465156 116164 465158
rect 116228 465156 116275 465160
rect 118510 465158 118556 465218
rect 118620 465216 118667 465220
rect 128670 465218 128676 465220
rect 118662 465160 118667 465216
rect 118550 465156 118556 465158
rect 118620 465156 118667 465160
rect 128630 465158 128676 465218
rect 128740 465216 128787 465220
rect 136030 465218 136036 465220
rect 128782 465160 128787 465216
rect 128670 465156 128676 465158
rect 128740 465156 128787 465160
rect 135990 465158 136036 465218
rect 136100 465216 136147 465220
rect 140998 465218 141004 465220
rect 136142 465160 136147 465216
rect 136030 465156 136036 465158
rect 136100 465156 136147 465160
rect 140958 465158 141004 465218
rect 141068 465216 141115 465220
rect 143574 465218 143580 465220
rect 141110 465160 141115 465216
rect 140998 465156 141004 465158
rect 141068 465156 141115 465160
rect 143534 465158 143580 465218
rect 143644 465216 143691 465220
rect 153326 465218 153332 465220
rect 143686 465160 143691 465216
rect 143574 465156 143580 465158
rect 143644 465156 143691 465160
rect 153286 465158 153332 465218
rect 153396 465216 153443 465220
rect 156086 465218 156092 465220
rect 153438 465160 153443 465216
rect 153326 465156 153332 465158
rect 153396 465156 153443 465160
rect 156046 465158 156092 465218
rect 156156 465216 156203 465220
rect 168414 465218 168420 465220
rect 156198 465160 156203 465216
rect 156086 465156 156092 465158
rect 156156 465156 156203 465160
rect 168374 465158 168420 465218
rect 168484 465216 168531 465220
rect 169702 465218 169708 465220
rect 168526 465160 168531 465216
rect 168414 465156 168420 465158
rect 168484 465156 168531 465160
rect 169662 465158 169708 465218
rect 169772 465216 169819 465220
rect 169814 465160 169819 465216
rect 169702 465156 169708 465158
rect 169772 465156 169819 465160
rect 180926 465156 180932 465220
rect 180996 465218 181002 465220
rect 187693 465218 187759 465221
rect 180996 465216 187759 465218
rect 180996 465160 187698 465216
rect 187754 465160 187759 465216
rect 180996 465158 187759 465160
rect 180996 465156 181002 465158
rect 103697 465155 103763 465156
rect 111057 465155 111123 465156
rect 113817 465155 113883 465156
rect 116209 465155 116275 465156
rect 118601 465155 118667 465156
rect 128721 465155 128787 465156
rect 136081 465155 136147 465156
rect 141049 465155 141115 465156
rect 143625 465155 143691 465156
rect 153377 465155 153443 465156
rect 156137 465155 156203 465156
rect 168465 465155 168531 465156
rect 169753 465155 169819 465156
rect 187693 465155 187759 465158
rect 131113 463996 131179 463997
rect 131062 463994 131068 463996
rect 131022 463934 131068 463994
rect 131132 463992 131179 463996
rect 131174 463936 131179 463992
rect 131062 463932 131068 463934
rect 131132 463932 131179 463936
rect 131113 463931 131179 463932
rect 83457 463724 83523 463725
rect 120993 463724 121059 463725
rect 123569 463724 123635 463725
rect 125961 463724 126027 463725
rect 133505 463724 133571 463725
rect 138473 463724 138539 463725
rect 146017 463724 146083 463725
rect 148501 463724 148567 463725
rect 151077 463724 151143 463725
rect 83456 463660 83462 463724
rect 83526 463722 83532 463724
rect 83526 463662 83614 463722
rect 83526 463660 83532 463662
rect 120992 463660 120998 463724
rect 121062 463722 121068 463724
rect 121062 463662 121150 463722
rect 123569 463720 123582 463724
rect 123646 463722 123652 463724
rect 125888 463722 125894 463724
rect 123569 463664 123574 463720
rect 121062 463660 121068 463662
rect 123569 463660 123582 463664
rect 123646 463662 123726 463722
rect 125870 463662 125894 463722
rect 123646 463660 123652 463662
rect 125888 463660 125894 463662
rect 125958 463720 126027 463724
rect 125958 463664 125966 463720
rect 126022 463664 126027 463720
rect 125958 463660 126027 463664
rect 133504 463660 133510 463724
rect 133574 463722 133580 463724
rect 138400 463722 138406 463724
rect 133574 463662 133662 463722
rect 138382 463662 138406 463722
rect 133574 463660 133580 463662
rect 138400 463660 138406 463662
rect 138470 463720 138539 463724
rect 138470 463664 138478 463720
rect 138534 463664 138539 463720
rect 138470 463660 138539 463664
rect 146016 463660 146022 463724
rect 146086 463722 146092 463724
rect 148464 463722 148470 463724
rect 146086 463662 146174 463722
rect 148410 463662 148470 463722
rect 148534 463720 148567 463724
rect 151048 463722 151054 463724
rect 148562 463664 148567 463720
rect 146086 463660 146092 463662
rect 148464 463660 148470 463662
rect 148534 463660 148567 463664
rect 150986 463662 151054 463722
rect 151118 463720 151143 463724
rect 151138 463664 151143 463720
rect 151048 463660 151054 463662
rect 151118 463660 151143 463664
rect 83457 463659 83523 463660
rect 120993 463659 121059 463660
rect 123569 463659 123635 463660
rect 125961 463659 126027 463660
rect 133505 463659 133571 463660
rect 138473 463659 138539 463660
rect 146017 463659 146083 463660
rect 148501 463659 148567 463660
rect 151077 463659 151143 463660
rect -960 462634 480 462724
rect 3693 462634 3759 462637
rect -960 462632 3759 462634
rect -960 462576 3698 462632
rect 3754 462576 3759 462632
rect -960 462574 3759 462576
rect -960 462484 480 462574
rect 3693 462571 3759 462574
rect 186865 461546 186931 461549
rect 238150 461546 238156 461548
rect 186865 461544 238156 461546
rect 186865 461488 186870 461544
rect 186926 461488 238156 461544
rect 186865 461486 238156 461488
rect 186865 461483 186931 461486
rect 238150 461484 238156 461486
rect 238220 461484 238226 461548
rect 189073 459234 189139 459237
rect 187190 459232 189139 459234
rect 187190 459220 189078 459232
rect 186588 459176 189078 459220
rect 189134 459176 189139 459232
rect 186588 459174 189139 459176
rect 186588 459160 187250 459174
rect 189073 459171 189139 459174
rect 583520 457996 584960 458236
rect -960 449578 480 449668
rect 2957 449578 3023 449581
rect -960 449576 3023 449578
rect -960 449520 2962 449576
rect 3018 449520 3023 449576
rect -960 449518 3023 449520
rect -960 449428 480 449518
rect 2957 449515 3023 449518
rect 583520 444668 584960 444908
rect 238569 440194 238635 440197
rect 238569 440192 240242 440194
rect 238569 440136 238574 440192
rect 238630 440136 240242 440192
rect 238569 440134 240242 440136
rect 238569 440131 238635 440134
rect 240182 439552 240242 440134
rect 237465 438154 237531 438157
rect 240182 438154 240242 438712
rect 237465 438152 240242 438154
rect 237465 438096 237470 438152
rect 237526 438096 240242 438152
rect 237465 438094 240242 438096
rect 237465 438091 237531 438094
rect 237373 437610 237439 437613
rect 240182 437610 240242 437760
rect 237373 437608 240242 437610
rect 237373 437552 237378 437608
rect 237434 437552 240242 437608
rect 237373 437550 240242 437552
rect 237373 437547 237439 437550
rect -960 436508 480 436748
rect 490414 435916 490420 435980
rect 490484 435978 490490 435980
rect 491518 435978 491524 435980
rect 490484 435918 491524 435978
rect 490484 435916 490490 435918
rect 491518 435916 491524 435918
rect 491588 435916 491594 435980
rect 238477 435842 238543 435845
rect 238477 435840 240242 435842
rect 238477 435784 238482 435840
rect 238538 435784 240242 435840
rect 238477 435782 240242 435784
rect 238477 435779 238543 435782
rect 240182 435232 240242 435782
rect 237465 433666 237531 433669
rect 240182 433666 240242 434224
rect 237465 433664 240242 433666
rect 237465 433608 237470 433664
rect 237526 433608 240242 433664
rect 237465 433606 240242 433608
rect 237465 433603 237531 433606
rect 237373 433394 237439 433397
rect 240182 433394 240242 433408
rect 237373 433392 240242 433394
rect 237373 433336 237378 433392
rect 237434 433336 240242 433392
rect 237373 433334 240242 433336
rect 237373 433331 237439 433334
rect 580901 431626 580967 431629
rect 583520 431626 584960 431716
rect 580901 431624 584960 431626
rect 580901 431568 580906 431624
rect 580962 431568 584960 431624
rect 580901 431566 584960 431568
rect 580901 431563 580967 431566
rect 583520 431476 584960 431566
rect 237373 431354 237439 431357
rect 237373 431352 240242 431354
rect 237373 431296 237378 431352
rect 237434 431296 240242 431352
rect 237373 431294 240242 431296
rect 237373 431291 237439 431294
rect 240182 430744 240242 431294
rect 237373 429314 237439 429317
rect 240182 429314 240242 429872
rect 237373 429312 240242 429314
rect 237373 429256 237378 429312
rect 237434 429256 240242 429312
rect 237373 429254 240242 429256
rect 237373 429251 237439 429254
rect 237373 428498 237439 428501
rect 240182 428498 240242 429056
rect 237373 428496 240242 428498
rect 237373 428440 237378 428496
rect 237434 428440 240242 428496
rect 237373 428438 240242 428440
rect 237373 428435 237439 428438
rect 237373 426322 237439 426325
rect 240182 426322 240242 426336
rect 237373 426320 240242 426322
rect 237373 426264 237378 426320
rect 237434 426264 240242 426320
rect 237373 426262 240242 426264
rect 237373 426259 237439 426262
rect 237373 425234 237439 425237
rect 240182 425234 240242 425520
rect 237373 425232 240242 425234
rect 237373 425176 237378 425232
rect 237434 425176 240242 425232
rect 237373 425174 240242 425176
rect 237373 425171 237439 425174
rect 237373 424010 237439 424013
rect 240182 424010 240242 424568
rect 237373 424008 240242 424010
rect 237373 423952 237378 424008
rect 237434 423952 240242 424008
rect 237373 423950 240242 423952
rect 237373 423947 237439 423950
rect -960 423452 480 423692
rect 237373 422106 237439 422109
rect 237373 422104 240242 422106
rect 237373 422048 237378 422104
rect 237434 422048 240242 422104
rect 237373 422046 240242 422048
rect 237373 422043 237439 422046
rect 240182 422040 240242 422046
rect 237373 421018 237439 421021
rect 240182 421018 240242 421032
rect 237373 421016 240242 421018
rect 237373 420960 237378 421016
rect 237434 420960 240242 421016
rect 237373 420958 240242 420960
rect 237373 420955 237439 420958
rect 237373 419658 237439 419661
rect 240182 419658 240242 420216
rect 237373 419656 240242 419658
rect 237373 419600 237378 419656
rect 237434 419600 240242 419656
rect 237373 419598 240242 419600
rect 237373 419595 237439 419598
rect 580165 418298 580231 418301
rect 583520 418298 584960 418388
rect 580165 418296 584960 418298
rect 580165 418240 580170 418296
rect 580226 418240 584960 418296
rect 580165 418238 584960 418240
rect 580165 418235 580231 418238
rect 238385 418162 238451 418165
rect 238385 418160 240242 418162
rect 238385 418104 238390 418160
rect 238446 418104 240242 418160
rect 583520 418148 584960 418238
rect 238385 418102 240242 418104
rect 238385 418099 238451 418102
rect 240182 417688 240242 418102
rect 48037 416938 48103 416941
rect 48037 416936 49434 416938
rect 48037 416880 48042 416936
rect 48098 416924 49434 416936
rect 48098 416880 50048 416924
rect 48037 416878 50048 416880
rect 48037 416875 48103 416878
rect 49374 416864 50048 416878
rect 237465 416122 237531 416125
rect 240182 416122 240242 416680
rect 237465 416120 240242 416122
rect 237465 416064 237470 416120
rect 237526 416064 240242 416120
rect 237465 416062 240242 416064
rect 237465 416059 237531 416062
rect 48129 415986 48195 415989
rect 48129 415984 49434 415986
rect 48129 415928 48134 415984
rect 48190 415972 49434 415984
rect 48190 415928 50048 415972
rect 48129 415926 50048 415928
rect 48129 415923 48195 415926
rect 49374 415912 50048 415926
rect 237373 415578 237439 415581
rect 240182 415578 240242 415864
rect 237373 415576 240242 415578
rect 237373 415520 237378 415576
rect 237434 415520 240242 415576
rect 237373 415518 240242 415520
rect 237373 415515 237439 415518
rect 47945 413810 48011 413813
rect 237373 413810 237439 413813
rect 47945 413808 49434 413810
rect 47945 413752 47950 413808
rect 48006 413796 49434 413808
rect 237373 413808 240242 413810
rect 48006 413752 50048 413796
rect 47945 413750 50048 413752
rect 47945 413747 48011 413750
rect 49374 413736 50048 413750
rect 237373 413752 237378 413808
rect 237434 413752 240242 413808
rect 237373 413750 240242 413752
rect 237373 413747 237439 413750
rect 240182 413200 240242 413750
rect 49325 412858 49391 412861
rect 49325 412856 49802 412858
rect 49325 412800 49330 412856
rect 49386 412844 49802 412856
rect 49386 412800 50048 412844
rect 49325 412798 50048 412800
rect 49325 412795 49391 412798
rect 49742 412784 50048 412798
rect 237373 411770 237439 411773
rect 240182 411770 240242 412328
rect 237373 411768 240242 411770
rect 237373 411712 237378 411768
rect 237434 411712 240242 411768
rect 237373 411710 240242 411712
rect 237373 411707 237439 411710
rect 238385 411362 238451 411365
rect 240182 411362 240242 411376
rect 238385 411360 240242 411362
rect 238385 411304 238390 411360
rect 238446 411304 240242 411360
rect 238385 411302 240242 411304
rect 238385 411299 238451 411302
rect 49417 411076 49483 411079
rect 49417 411074 50048 411076
rect 49417 411018 49422 411074
rect 49478 411018 50048 411074
rect 49417 411016 50048 411018
rect 49417 411013 49483 411016
rect -960 410546 480 410636
rect 3877 410546 3943 410549
rect -960 410544 3943 410546
rect -960 410488 3882 410544
rect 3938 410488 3943 410544
rect -960 410486 3943 410488
rect -960 410396 480 410486
rect 3877 410483 3943 410486
rect 49233 410002 49299 410005
rect 49233 410000 49802 410002
rect 49233 409944 49238 410000
rect 49294 409988 49802 410000
rect 49294 409944 50048 409988
rect 49233 409942 50048 409944
rect 49233 409939 49299 409942
rect 49742 409928 50048 409942
rect 238293 409458 238359 409461
rect 238293 409456 240242 409458
rect 238293 409400 238298 409456
rect 238354 409400 240242 409456
rect 238293 409398 240242 409400
rect 238293 409395 238359 409398
rect 240182 408848 240242 409398
rect 49601 408220 49667 408223
rect 49601 408218 50048 408220
rect 49601 408162 49606 408218
rect 49662 408162 50048 408218
rect 49601 408160 50048 408162
rect 49601 408157 49667 408160
rect 237373 407418 237439 407421
rect 240182 407418 240242 407976
rect 237373 407416 240242 407418
rect 237373 407360 237378 407416
rect 237434 407360 240242 407416
rect 237373 407358 240242 407360
rect 237373 407355 237439 407358
rect 238293 406466 238359 406469
rect 240182 406466 240242 407024
rect 238293 406464 240242 406466
rect 238293 406408 238298 406464
rect 238354 406408 240242 406464
rect 238293 406406 240242 406408
rect 238293 406403 238359 406406
rect 237373 405106 237439 405109
rect 237373 405104 240242 405106
rect 237373 405048 237378 405104
rect 237434 405048 240242 405104
rect 237373 405046 240242 405048
rect 237373 405043 237439 405046
rect 240182 404496 240242 405046
rect 583520 404820 584960 405060
rect 237373 403338 237439 403341
rect 240182 403338 240242 403488
rect 237373 403336 240242 403338
rect 237373 403280 237378 403336
rect 237434 403280 240242 403336
rect 237373 403278 240242 403280
rect 237373 403275 237439 403278
rect 238477 402114 238543 402117
rect 240182 402114 240242 402672
rect 238477 402112 240242 402114
rect 238477 402056 238482 402112
rect 238538 402056 240242 402112
rect 238477 402054 240242 402056
rect 238477 402051 238543 402054
rect 237373 400074 237439 400077
rect 237373 400072 240242 400074
rect 237373 400016 237378 400072
rect 237434 400016 240242 400072
rect 237373 400014 240242 400016
rect 237373 400011 237439 400014
rect 240182 400008 240242 400014
rect 189073 399394 189139 399397
rect 187190 399392 189139 399394
rect 187190 399380 189078 399392
rect 186588 399336 189078 399380
rect 189134 399336 189139 399392
rect 186588 399334 189139 399336
rect 186588 399320 187250 399334
rect 189073 399331 189139 399334
rect 237373 398986 237439 398989
rect 240182 398986 240242 399136
rect 237373 398984 240242 398986
rect 237373 398928 237378 398984
rect 237434 398928 240242 398984
rect 237373 398926 240242 398928
rect 237373 398923 237439 398926
rect 189073 397762 189139 397765
rect 187190 397760 189139 397762
rect 187190 397748 189078 397760
rect 186588 397704 189078 397748
rect 189134 397704 189139 397760
rect 186588 397702 189139 397704
rect 186588 397688 187250 397702
rect 189073 397699 189139 397702
rect 238569 397626 238635 397629
rect 240182 397626 240242 398184
rect 238569 397624 240242 397626
rect -960 397490 480 397580
rect 238569 397568 238574 397624
rect 238630 397568 240242 397624
rect 238569 397566 240242 397568
rect 238569 397563 238635 397566
rect 3325 397490 3391 397493
rect -960 397488 3391 397490
rect -960 397432 3330 397488
rect 3386 397432 3391 397488
rect -960 397430 3391 397432
rect -960 397340 480 397430
rect 3325 397427 3391 397430
rect 189257 396402 189323 396405
rect 187190 396400 189323 396402
rect 187190 396388 189262 396400
rect 186588 396344 189262 396388
rect 189318 396344 189323 396400
rect 186588 396342 189323 396344
rect 186588 396328 187250 396342
rect 189257 396339 189323 396342
rect 237373 395994 237439 395997
rect 237373 395992 240242 395994
rect 237373 395936 237378 395992
rect 237434 395936 240242 395992
rect 237373 395934 240242 395936
rect 237373 395931 237439 395934
rect 240182 395656 240242 395934
rect 189073 394906 189139 394909
rect 187190 394904 189139 394906
rect 187190 394892 189078 394904
rect 186588 394848 189078 394892
rect 189134 394848 189139 394904
rect 186588 394846 189139 394848
rect 186588 394832 187250 394846
rect 189073 394843 189139 394846
rect 237373 394770 237439 394773
rect 240182 394770 240242 394784
rect 237373 394768 240242 394770
rect 237373 394712 237378 394768
rect 237434 394712 240242 394768
rect 237373 394710 240242 394712
rect 237373 394707 237439 394710
rect 189257 393682 189323 393685
rect 187190 393680 189323 393682
rect 187190 393668 189262 393680
rect 186588 393624 189262 393668
rect 189318 393624 189323 393680
rect 186588 393622 189323 393624
rect 186588 393608 187250 393622
rect 189257 393619 189323 393622
rect 238661 393410 238727 393413
rect 240182 393410 240242 393832
rect 238661 393408 240242 393410
rect 238661 393352 238666 393408
rect 238722 393352 240242 393408
rect 238661 393350 240242 393352
rect 238661 393347 238727 393350
rect 237373 391914 237439 391917
rect 237373 391912 240242 391914
rect 237373 391856 237378 391912
rect 237434 391856 240242 391912
rect 237373 391854 240242 391856
rect 237373 391851 237439 391854
rect 240182 391304 240242 391854
rect 583520 391628 584960 391868
rect 48221 390010 48287 390013
rect 48221 390008 49434 390010
rect 48221 389952 48226 390008
rect 48282 389996 49434 390008
rect 48282 389952 50048 389996
rect 48221 389950 50048 389952
rect 48221 389947 48287 389950
rect 49374 389936 50048 389950
rect 237465 389738 237531 389741
rect 240182 389738 240242 390296
rect 237465 389736 240242 389738
rect 237465 389680 237470 389736
rect 237526 389680 240242 389736
rect 237465 389678 240242 389680
rect 237465 389675 237531 389678
rect 237373 389330 237439 389333
rect 240182 389330 240242 389480
rect 237373 389328 240242 389330
rect 237373 389272 237378 389328
rect 237434 389272 240242 389328
rect 237373 389270 240242 389272
rect 237373 389267 237439 389270
rect 47577 388378 47643 388381
rect 47577 388376 49434 388378
rect 47577 388320 47582 388376
rect 47638 388364 49434 388376
rect 47638 388320 50048 388364
rect 47577 388318 50048 388320
rect 47577 388315 47643 388318
rect 49374 388304 50048 388318
rect 47853 388106 47919 388109
rect 47853 388104 49434 388106
rect 47853 388048 47858 388104
rect 47914 388092 49434 388104
rect 47914 388048 50048 388092
rect 47853 388046 50048 388048
rect 47853 388043 47919 388046
rect 49374 388032 50048 388046
rect 237373 387426 237439 387429
rect 237373 387424 240242 387426
rect 237373 387368 237378 387424
rect 237434 387368 240242 387424
rect 237373 387366 240242 387368
rect 237373 387363 237439 387366
rect 240182 386816 240242 387366
rect 237373 385386 237439 385389
rect 240182 385386 240242 385944
rect 237373 385384 240242 385386
rect 237373 385328 237378 385384
rect 237434 385328 240242 385384
rect 237373 385326 240242 385328
rect 237373 385323 237439 385326
rect 237465 385114 237531 385117
rect 240182 385114 240242 385128
rect 237465 385112 240242 385114
rect 237465 385056 237470 385112
rect 237526 385056 240242 385112
rect 237465 385054 240242 385056
rect 237465 385051 237531 385054
rect -960 384284 480 384524
rect 237373 383074 237439 383077
rect 237373 383072 240242 383074
rect 237373 383016 237378 383072
rect 237434 383016 240242 383072
rect 237373 383014 240242 383016
rect 237373 383011 237439 383014
rect 240182 382464 240242 383014
rect 237373 381034 237439 381037
rect 240182 381034 240242 381592
rect 237373 381032 240242 381034
rect 237373 380976 237378 381032
rect 237434 380976 240242 381032
rect 237373 380974 240242 380976
rect 237373 380971 237439 380974
rect 237373 380082 237439 380085
rect 240182 380082 240242 380640
rect 237373 380080 240242 380082
rect 237373 380024 237378 380080
rect 237434 380024 240242 380080
rect 237373 380022 240242 380024
rect 237373 380019 237439 380022
rect 123477 379676 123543 379677
rect 130929 379676 130995 379677
rect 133505 379676 133571 379677
rect 145925 379676 145991 379677
rect 148501 379676 148567 379677
rect 155953 379676 156019 379677
rect 123440 379674 123446 379676
rect 123386 379614 123446 379674
rect 123510 379672 123543 379676
rect 130920 379674 130926 379676
rect 123538 379616 123543 379672
rect 123440 379612 123446 379614
rect 123510 379612 123543 379616
rect 130838 379614 130926 379674
rect 130920 379612 130926 379614
rect 130990 379612 130996 379676
rect 133504 379612 133510 379676
rect 133574 379674 133580 379676
rect 145880 379674 145886 379676
rect 133574 379614 133662 379674
rect 145834 379614 145886 379674
rect 145950 379672 145991 379676
rect 148464 379674 148470 379676
rect 145986 379616 145991 379672
rect 133574 379612 133580 379614
rect 145880 379612 145886 379614
rect 145950 379612 145991 379616
rect 148410 379614 148470 379674
rect 148534 379672 148567 379676
rect 155944 379674 155950 379676
rect 148562 379616 148567 379672
rect 148464 379612 148470 379614
rect 148534 379612 148567 379616
rect 155862 379614 155950 379674
rect 155944 379612 155950 379614
rect 156014 379612 156020 379676
rect 123477 379611 123543 379612
rect 130929 379611 130995 379612
rect 133505 379611 133571 379612
rect 145925 379611 145991 379612
rect 148501 379611 148567 379612
rect 155953 379611 156019 379612
rect 93945 379540 94011 379541
rect 96429 379540 96495 379541
rect 97625 379540 97691 379541
rect 98729 379540 98795 379541
rect 102225 379540 102291 379541
rect 125961 379540 126027 379541
rect 128537 379540 128603 379541
rect 93928 379538 93934 379540
rect 93854 379478 93934 379538
rect 93998 379536 94011 379540
rect 96376 379538 96382 379540
rect 94006 379480 94011 379536
rect 93928 379476 93934 379478
rect 93998 379476 94011 379480
rect 96338 379478 96382 379538
rect 96446 379536 96495 379540
rect 97600 379538 97606 379540
rect 96490 379480 96495 379536
rect 96376 379476 96382 379478
rect 96446 379476 96495 379480
rect 97534 379478 97606 379538
rect 97670 379536 97691 379540
rect 98688 379538 98694 379540
rect 97686 379480 97691 379536
rect 97600 379476 97606 379478
rect 97670 379476 97691 379480
rect 98638 379478 98694 379538
rect 98758 379536 98795 379540
rect 98790 379480 98795 379536
rect 98688 379476 98694 379478
rect 98758 379476 98795 379480
rect 102224 379476 102230 379540
rect 102294 379538 102300 379540
rect 125910 379538 125916 379540
rect 102294 379478 102382 379538
rect 125870 379478 125916 379538
rect 125980 379536 126027 379540
rect 128486 379538 128492 379540
rect 126022 379480 126027 379536
rect 102294 379476 102300 379478
rect 125910 379476 125916 379478
rect 125980 379476 126027 379480
rect 128446 379478 128492 379538
rect 128556 379536 128603 379540
rect 128598 379480 128603 379536
rect 128486 379476 128492 379478
rect 128556 379476 128603 379480
rect 93945 379475 94011 379476
rect 96429 379475 96495 379476
rect 97625 379475 97691 379476
rect 98729 379475 98795 379476
rect 102225 379475 102291 379476
rect 125961 379475 126027 379476
rect 128537 379475 128603 379476
rect 108062 379340 108068 379404
rect 108132 379402 108138 379404
rect 191189 379402 191255 379405
rect 108132 379400 191255 379402
rect 108132 379344 191194 379400
rect 191250 379344 191255 379400
rect 108132 379342 191255 379344
rect 108132 379340 108138 379342
rect 191189 379339 191255 379342
rect 150985 379268 151051 379269
rect 150934 379266 150940 379268
rect 150894 379206 150940 379266
rect 151004 379264 151051 379268
rect 151046 379208 151051 379264
rect 150934 379204 150940 379206
rect 151004 379204 151051 379208
rect 150985 379203 151051 379204
rect 579797 378450 579863 378453
rect 583520 378450 584960 378540
rect 579797 378448 584960 378450
rect 579797 378392 579802 378448
rect 579858 378392 584960 378448
rect 579797 378390 584960 378392
rect 579797 378387 579863 378390
rect 583520 378300 584960 378390
rect 67214 378116 67220 378180
rect 67284 378116 67290 378180
rect 74206 378116 74212 378180
rect 74276 378116 74282 378180
rect 77702 378116 77708 378180
rect 77772 378116 77778 378180
rect 81198 378116 81204 378180
rect 81268 378116 81274 378180
rect 91870 378116 91876 378180
rect 91940 378116 91946 378180
rect 95918 378116 95924 378180
rect 95988 378116 95994 378180
rect 99782 378116 99788 378180
rect 99852 378116 99858 378180
rect 103278 378116 103284 378180
rect 103348 378116 103354 378180
rect 103646 378116 103652 378180
rect 103716 378116 103722 378180
rect 113582 378116 113588 378180
rect 113652 378116 113658 378180
rect 120942 378116 120948 378180
rect 121012 378116 121018 378180
rect 153326 378116 153332 378180
rect 153396 378116 153402 378180
rect 67222 378042 67282 378116
rect 67541 378042 67607 378045
rect 73153 378044 73219 378045
rect 73102 378042 73108 378044
rect 67222 378040 67607 378042
rect 67222 377984 67546 378040
rect 67602 377984 67607 378040
rect 67222 377982 67607 377984
rect 73062 377982 73108 378042
rect 73172 378040 73219 378044
rect 73214 377984 73219 378040
rect 67541 377979 67607 377982
rect 73102 377980 73108 377982
rect 73172 377980 73219 377984
rect 74214 378042 74274 378116
rect 74349 378042 74415 378045
rect 74214 378040 74415 378042
rect 74214 377984 74354 378040
rect 74410 377984 74415 378040
rect 74214 377982 74415 377984
rect 77710 378042 77770 378116
rect 81206 378045 81266 378116
rect 78489 378042 78555 378045
rect 77710 378040 78555 378042
rect 77710 377984 78494 378040
rect 78550 377984 78555 378040
rect 77710 377982 78555 377984
rect 73153 377979 73219 377980
rect 74349 377979 74415 377982
rect 78489 377979 78555 377982
rect 81157 378040 81266 378045
rect 81157 377984 81162 378040
rect 81218 377984 81266 378040
rect 81157 377982 81266 377984
rect 91878 378042 91938 378116
rect 92289 378042 92355 378045
rect 92841 378044 92907 378045
rect 92790 378042 92796 378044
rect 91878 378040 92355 378042
rect 91878 377984 92294 378040
rect 92350 377984 92355 378040
rect 91878 377982 92355 377984
rect 92750 377982 92796 378042
rect 92860 378040 92907 378044
rect 92902 377984 92907 378040
rect 81157 377979 81223 377982
rect 92289 377979 92355 377982
rect 92790 377980 92796 377982
rect 92860 377980 92907 377984
rect 95182 377980 95188 378044
rect 95252 378042 95258 378044
rect 95325 378042 95391 378045
rect 95252 378040 95391 378042
rect 95252 377984 95330 378040
rect 95386 377984 95391 378040
rect 95252 377982 95391 377984
rect 95926 378042 95986 378116
rect 99790 378045 99850 378116
rect 103286 378045 103346 378116
rect 96521 378042 96587 378045
rect 95926 378040 96587 378042
rect 95926 377984 96526 378040
rect 96582 377984 96587 378040
rect 95926 377982 96587 377984
rect 99790 378040 99899 378045
rect 101305 378044 101371 378045
rect 101254 378042 101260 378044
rect 99790 377984 99838 378040
rect 99894 377984 99899 378040
rect 99790 377982 99899 377984
rect 101214 377982 101260 378042
rect 101324 378040 101371 378044
rect 101366 377984 101371 378040
rect 95252 377980 95258 377982
rect 92841 377979 92907 377980
rect 95325 377979 95391 377982
rect 96521 377979 96587 377982
rect 99833 377979 99899 377982
rect 101254 377980 101260 377982
rect 101324 377980 101371 377984
rect 103286 378040 103395 378045
rect 103286 377984 103334 378040
rect 103390 377984 103395 378040
rect 103286 377982 103395 377984
rect 103654 378042 103714 378116
rect 104801 378042 104867 378045
rect 105905 378044 105971 378045
rect 105854 378042 105860 378044
rect 103654 378040 104867 378042
rect 103654 377984 104806 378040
rect 104862 377984 104867 378040
rect 103654 377982 104867 377984
rect 105814 377982 105860 378042
rect 105924 378040 105971 378044
rect 105966 377984 105971 378040
rect 101305 377979 101371 377980
rect 103329 377979 103395 377982
rect 104801 377979 104867 377982
rect 105854 377980 105860 377982
rect 105924 377980 105971 377984
rect 106958 377980 106964 378044
rect 107028 378042 107034 378044
rect 107561 378042 107627 378045
rect 107028 378040 107627 378042
rect 107028 377984 107566 378040
rect 107622 377984 107627 378040
rect 107028 377982 107627 377984
rect 107028 377980 107034 377982
rect 105905 377979 105971 377980
rect 107561 377979 107627 377982
rect 109166 377980 109172 378044
rect 109236 378042 109242 378044
rect 110229 378042 110295 378045
rect 109236 378040 110295 378042
rect 109236 377984 110234 378040
rect 110290 377984 110295 378040
rect 109236 377982 110295 377984
rect 113590 378042 113650 378116
rect 120950 378045 121010 378116
rect 153334 378045 153394 378116
rect 114461 378042 114527 378045
rect 113590 378040 114527 378042
rect 113590 377984 114466 378040
rect 114522 377984 114527 378040
rect 113590 377982 114527 377984
rect 120950 378040 121059 378045
rect 136081 378044 136147 378045
rect 136030 378042 136036 378044
rect 120950 377984 120998 378040
rect 121054 377984 121059 378040
rect 120950 377982 121059 377984
rect 135990 377982 136036 378042
rect 136100 378040 136147 378044
rect 136142 377984 136147 378040
rect 109236 377980 109242 377982
rect 110229 377979 110295 377982
rect 114461 377979 114527 377982
rect 120993 377979 121059 377982
rect 136030 377980 136036 377982
rect 136100 377980 136147 377984
rect 138606 377980 138612 378044
rect 138676 378042 138682 378044
rect 139025 378042 139091 378045
rect 138676 378040 139091 378042
rect 138676 377984 139030 378040
rect 139086 377984 139091 378040
rect 138676 377982 139091 377984
rect 138676 377980 138682 377982
rect 136081 377979 136147 377980
rect 139025 377979 139091 377982
rect 140998 377980 141004 378044
rect 141068 378042 141074 378044
rect 141601 378042 141667 378045
rect 143441 378044 143507 378045
rect 143390 378042 143396 378044
rect 141068 378040 141667 378042
rect 141068 377984 141606 378040
rect 141662 377984 141667 378040
rect 141068 377982 141667 377984
rect 143350 377982 143396 378042
rect 143460 378040 143507 378044
rect 143502 377984 143507 378040
rect 141068 377980 141074 377982
rect 141601 377979 141667 377982
rect 143390 377980 143396 377982
rect 143460 377980 143507 377984
rect 153334 378040 153443 378045
rect 153334 377984 153382 378040
rect 153438 377984 153443 378040
rect 153334 377982 153443 377984
rect 143441 377979 143507 377980
rect 153377 377979 153443 377982
rect 104433 377908 104499 377909
rect 104382 377906 104388 377908
rect 104342 377846 104388 377906
rect 104452 377904 104499 377908
rect 104494 377848 104499 377904
rect 104382 377844 104388 377846
rect 104452 377844 104499 377848
rect 104433 377843 104499 377844
rect 240182 377498 240242 378056
rect 219390 377438 240242 377498
rect 180701 377362 180767 377365
rect 187693 377362 187759 377365
rect 180701 377360 187759 377362
rect 180701 377304 180706 377360
rect 180762 377304 187698 377360
rect 187754 377304 187759 377360
rect 180701 377302 187759 377304
rect 180701 377299 180767 377302
rect 187693 377299 187759 377302
rect 66161 377092 66227 377093
rect 66110 377090 66116 377092
rect 66070 377030 66116 377090
rect 66180 377088 66227 377092
rect 66222 377032 66227 377088
rect 66110 377028 66116 377030
rect 66180 377028 66227 377032
rect 68318 377028 68324 377092
rect 68388 377090 68394 377092
rect 68921 377090 68987 377093
rect 68388 377088 68987 377090
rect 68388 377032 68926 377088
rect 68982 377032 68987 377088
rect 68388 377030 68987 377032
rect 68388 377028 68394 377030
rect 66161 377027 66227 377028
rect 68921 377027 68987 377030
rect 69606 377028 69612 377092
rect 69676 377090 69682 377092
rect 70301 377090 70367 377093
rect 69676 377088 70367 377090
rect 69676 377032 70306 377088
rect 70362 377032 70367 377088
rect 69676 377030 70367 377032
rect 69676 377028 69682 377030
rect 70301 377027 70367 377030
rect 70526 377028 70532 377092
rect 70596 377090 70602 377092
rect 71681 377090 71747 377093
rect 70596 377088 71747 377090
rect 70596 377032 71686 377088
rect 71742 377032 71747 377088
rect 70596 377030 71747 377032
rect 70596 377028 70602 377030
rect 71681 377027 71747 377030
rect 71814 377028 71820 377092
rect 71884 377090 71890 377092
rect 73061 377090 73127 377093
rect 71884 377088 73127 377090
rect 71884 377032 73066 377088
rect 73122 377032 73127 377088
rect 71884 377030 73127 377032
rect 71884 377028 71890 377030
rect 73061 377027 73127 377030
rect 75494 377028 75500 377092
rect 75564 377090 75570 377092
rect 75821 377090 75887 377093
rect 75564 377088 75887 377090
rect 75564 377032 75826 377088
rect 75882 377032 75887 377088
rect 75564 377030 75887 377032
rect 75564 377028 75570 377030
rect 75821 377027 75887 377030
rect 76598 377028 76604 377092
rect 76668 377090 76674 377092
rect 77201 377090 77267 377093
rect 78305 377092 78371 377093
rect 78254 377090 78260 377092
rect 76668 377088 77267 377090
rect 76668 377032 77206 377088
rect 77262 377032 77267 377088
rect 76668 377030 77267 377032
rect 78214 377030 78260 377090
rect 78324 377088 78371 377092
rect 78366 377032 78371 377088
rect 76668 377028 76674 377030
rect 77201 377027 77267 377030
rect 78254 377028 78260 377030
rect 78324 377028 78371 377032
rect 78806 377028 78812 377092
rect 78876 377090 78882 377092
rect 79961 377090 80027 377093
rect 78876 377088 80027 377090
rect 78876 377032 79966 377088
rect 80022 377032 80027 377088
rect 78876 377030 80027 377032
rect 78876 377028 78882 377030
rect 78305 377027 78371 377028
rect 79961 377027 80027 377030
rect 80094 377028 80100 377092
rect 80164 377090 80170 377092
rect 81249 377090 81315 377093
rect 80164 377088 81315 377090
rect 80164 377032 81254 377088
rect 81310 377032 81315 377088
rect 80164 377030 81315 377032
rect 80164 377028 80170 377030
rect 81249 377027 81315 377030
rect 82486 377028 82492 377092
rect 82556 377090 82562 377092
rect 82721 377090 82787 377093
rect 82556 377088 82787 377090
rect 82556 377032 82726 377088
rect 82782 377032 82787 377088
rect 82556 377030 82787 377032
rect 82556 377028 82562 377030
rect 82721 377027 82787 377030
rect 83590 377028 83596 377092
rect 83660 377090 83666 377092
rect 84101 377090 84167 377093
rect 83660 377088 84167 377090
rect 83660 377032 84106 377088
rect 84162 377032 84167 377088
rect 83660 377030 84167 377032
rect 83660 377028 83666 377030
rect 84101 377027 84167 377030
rect 84510 377028 84516 377092
rect 84580 377090 84586 377092
rect 85481 377090 85547 377093
rect 84580 377088 85547 377090
rect 84580 377032 85486 377088
rect 85542 377032 85547 377088
rect 84580 377030 85547 377032
rect 84580 377028 84586 377030
rect 85481 377027 85547 377030
rect 85982 377028 85988 377092
rect 86052 377090 86058 377092
rect 86861 377090 86927 377093
rect 86052 377088 86927 377090
rect 86052 377032 86866 377088
rect 86922 377032 86927 377088
rect 86052 377030 86927 377032
rect 86052 377028 86058 377030
rect 86861 377027 86927 377030
rect 88006 377028 88012 377092
rect 88076 377090 88082 377092
rect 88149 377090 88215 377093
rect 89529 377092 89595 377093
rect 89478 377090 89484 377092
rect 88076 377088 88215 377090
rect 88076 377032 88154 377088
rect 88210 377032 88215 377088
rect 88076 377030 88215 377032
rect 89438 377030 89484 377090
rect 89548 377088 89595 377092
rect 89590 377032 89595 377088
rect 88076 377028 88082 377030
rect 88149 377027 88215 377030
rect 89478 377028 89484 377030
rect 89548 377028 89595 377032
rect 90766 377028 90772 377092
rect 90836 377090 90842 377092
rect 91001 377090 91067 377093
rect 90836 377088 91067 377090
rect 90836 377032 91006 377088
rect 91062 377032 91067 377088
rect 90836 377030 91067 377032
rect 90836 377028 90842 377030
rect 89529 377027 89595 377028
rect 91001 377027 91067 377030
rect 91134 377028 91140 377092
rect 91204 377090 91210 377092
rect 91737 377090 91803 377093
rect 91204 377088 91803 377090
rect 91204 377032 91742 377088
rect 91798 377032 91803 377088
rect 91204 377030 91803 377032
rect 91204 377028 91210 377030
rect 91737 377027 91803 377030
rect 93526 377028 93532 377092
rect 93596 377090 93602 377092
rect 93761 377090 93827 377093
rect 93596 377088 93827 377090
rect 93596 377032 93766 377088
rect 93822 377032 93827 377088
rect 93596 377030 93827 377032
rect 93596 377028 93602 377030
rect 93761 377027 93827 377030
rect 98310 377028 98316 377092
rect 98380 377090 98386 377092
rect 99281 377090 99347 377093
rect 98380 377088 99347 377090
rect 98380 377032 99286 377088
rect 99342 377032 99347 377088
rect 98380 377030 99347 377032
rect 98380 377028 98386 377030
rect 99281 377027 99347 377030
rect 101070 377028 101076 377092
rect 101140 377090 101146 377092
rect 102041 377090 102107 377093
rect 101140 377088 102107 377090
rect 101140 377032 102046 377088
rect 102102 377032 102107 377088
rect 101140 377030 102107 377032
rect 101140 377028 101146 377030
rect 102041 377027 102107 377030
rect 106038 377028 106044 377092
rect 106108 377090 106114 377092
rect 106181 377090 106247 377093
rect 106108 377088 106247 377090
rect 106108 377032 106186 377088
rect 106242 377032 106247 377088
rect 106108 377030 106247 377032
rect 106108 377028 106114 377030
rect 106181 377027 106247 377030
rect 108430 377028 108436 377092
rect 108500 377090 108506 377092
rect 108941 377090 109007 377093
rect 108500 377088 109007 377090
rect 108500 377032 108946 377088
rect 109002 377032 109007 377088
rect 108500 377030 109007 377032
rect 108500 377028 108506 377030
rect 108941 377027 109007 377030
rect 111006 377028 111012 377092
rect 111076 377090 111082 377092
rect 111701 377090 111767 377093
rect 111076 377088 111767 377090
rect 111076 377032 111706 377088
rect 111762 377032 111767 377088
rect 111076 377030 111767 377032
rect 111076 377028 111082 377030
rect 111701 377027 111767 377030
rect 115974 377028 115980 377092
rect 116044 377090 116050 377092
rect 117221 377090 117287 377093
rect 116044 377088 117287 377090
rect 116044 377032 117226 377088
rect 117282 377032 117287 377088
rect 116044 377030 117287 377032
rect 116044 377028 116050 377030
rect 117221 377027 117287 377030
rect 118366 377028 118372 377092
rect 118436 377090 118442 377092
rect 118601 377090 118667 377093
rect 118436 377088 118667 377090
rect 118436 377032 118606 377088
rect 118662 377032 118667 377088
rect 118436 377030 118667 377032
rect 118436 377028 118442 377030
rect 118601 377027 118667 377030
rect 173382 377028 173388 377092
rect 173452 377090 173458 377092
rect 173709 377090 173775 377093
rect 173452 377088 173775 377090
rect 173452 377032 173714 377088
rect 173770 377032 173775 377088
rect 173452 377030 173775 377032
rect 173452 377028 173458 377030
rect 173709 377027 173775 377030
rect 80830 376892 80836 376956
rect 80900 376954 80906 376956
rect 81341 376954 81407 376957
rect 80900 376952 81407 376954
rect 80900 376896 81346 376952
rect 81402 376896 81407 376952
rect 80900 376894 81407 376896
rect 80900 376892 80906 376894
rect 81341 376891 81407 376894
rect 83406 376892 83412 376956
rect 83476 376954 83482 376956
rect 84009 376954 84075 376957
rect 83476 376952 84075 376954
rect 83476 376896 84014 376952
rect 84070 376896 84075 376952
rect 83476 376894 84075 376896
rect 83476 376892 83482 376894
rect 84009 376891 84075 376894
rect 85798 376892 85804 376956
rect 85868 376954 85874 376956
rect 86769 376954 86835 376957
rect 85868 376952 86835 376954
rect 85868 376896 86774 376952
rect 86830 376896 86835 376952
rect 85868 376894 86835 376896
rect 85868 376892 85874 376894
rect 86769 376891 86835 376894
rect 87086 376892 87092 376956
rect 87156 376954 87162 376956
rect 88241 376954 88307 376957
rect 87156 376952 88307 376954
rect 87156 376896 88246 376952
rect 88302 376896 88307 376952
rect 87156 376894 88307 376896
rect 87156 376892 87162 376894
rect 88241 376891 88307 376894
rect 88558 376892 88564 376956
rect 88628 376954 88634 376956
rect 89621 376954 89687 376957
rect 88628 376952 89687 376954
rect 88628 376896 89626 376952
rect 89682 376896 89687 376952
rect 88628 376894 89687 376896
rect 88628 376892 88634 376894
rect 89621 376891 89687 376894
rect 173198 376892 173204 376956
rect 173268 376954 173274 376956
rect 173801 376954 173867 376957
rect 173268 376952 173867 376954
rect 173268 376896 173806 376952
rect 173862 376896 173867 376952
rect 173268 376894 173867 376896
rect 173268 376892 173274 376894
rect 173801 376891 173867 376894
rect 186957 376954 187023 376957
rect 219390 376954 219450 377438
rect 237373 377362 237439 377365
rect 237373 377360 240242 377362
rect 237373 377304 237378 377360
rect 237434 377304 240242 377360
rect 237373 377302 240242 377304
rect 237373 377299 237439 377302
rect 240182 377160 240242 377302
rect 186957 376952 219450 376954
rect 186957 376896 186962 376952
rect 187018 376896 219450 376952
rect 186957 376894 219450 376896
rect 186957 376891 187023 376894
rect 237373 376682 237439 376685
rect 237373 376680 240242 376682
rect 237373 376624 237378 376680
rect 237434 376624 240242 376680
rect 237373 376622 240242 376624
rect 237373 376619 237439 376622
rect 240182 376344 240242 376622
rect 238201 373962 238267 373965
rect 238201 373960 240242 373962
rect 238201 373904 238206 373960
rect 238262 373904 240242 373960
rect 238201 373902 240242 373904
rect 238201 373899 238267 373902
rect 240182 373760 240242 373902
rect 237373 373418 237439 373421
rect 237373 373416 240242 373418
rect 237373 373360 237378 373416
rect 237434 373360 240242 373416
rect 237373 373358 240242 373360
rect 237373 373355 237439 373358
rect 240182 372808 240242 373358
rect 237373 372330 237439 372333
rect 237373 372328 240242 372330
rect 237373 372272 237378 372328
rect 237434 372272 240242 372328
rect 237373 372270 240242 372272
rect 237373 372267 237439 372270
rect 240182 371992 240242 372270
rect -960 371228 480 371468
rect 238109 369746 238175 369749
rect 238109 369744 240242 369746
rect 238109 369688 238114 369744
rect 238170 369688 240242 369744
rect 238109 369686 240242 369688
rect 238109 369683 238175 369686
rect 240182 369272 240242 369686
rect 237373 368386 237439 368389
rect 240182 368386 240242 368400
rect 237373 368384 240242 368386
rect 237373 368328 237378 368384
rect 237434 368328 240242 368384
rect 237373 368326 240242 368328
rect 237373 368323 237439 368326
rect 237465 368114 237531 368117
rect 237465 368112 240242 368114
rect 237465 368056 237470 368112
rect 237526 368056 240242 368112
rect 237465 368054 240242 368056
rect 237465 368051 237531 368054
rect 240182 367504 240242 368054
rect 238017 365530 238083 365533
rect 238017 365528 240242 365530
rect 238017 365472 238022 365528
rect 238078 365472 240242 365528
rect 238017 365470 240242 365472
rect 238017 365467 238083 365470
rect 240182 364920 240242 365470
rect 580165 365122 580231 365125
rect 583520 365122 584960 365212
rect 580165 365120 584960 365122
rect 580165 365064 580170 365120
rect 580226 365064 584960 365120
rect 580165 365062 584960 365064
rect 580165 365059 580231 365062
rect 583520 364972 584960 365062
rect 237373 364170 237439 364173
rect 237373 364168 240242 364170
rect 237373 364112 237378 364168
rect 237434 364112 240242 364168
rect 237373 364110 240242 364112
rect 237373 364107 237439 364110
rect 240182 364104 240242 364110
rect 237465 363762 237531 363765
rect 237465 363760 240242 363762
rect 237465 363704 237470 363760
rect 237526 363704 240242 363760
rect 237465 363702 240242 363704
rect 237465 363699 237531 363702
rect 240182 363152 240242 363702
rect 237373 361178 237439 361181
rect 237373 361176 240242 361178
rect 237373 361120 237378 361176
rect 237434 361120 240242 361176
rect 237373 361118 240242 361120
rect 237373 361115 237439 361118
rect 240182 360568 240242 361118
rect 237373 359954 237439 359957
rect 237373 359952 240242 359954
rect 237373 359896 237378 359952
rect 237434 359896 240242 359952
rect 237373 359894 240242 359896
rect 237373 359891 237439 359894
rect 240182 359616 240242 359894
rect 237373 358730 237439 358733
rect 240182 358730 240242 358744
rect 237373 358728 240242 358730
rect 237373 358672 237378 358728
rect 237434 358672 240242 358728
rect 237373 358670 240242 358672
rect 237373 358667 237439 358670
rect -960 358458 480 358548
rect 3785 358458 3851 358461
rect -960 358456 3851 358458
rect -960 358400 3790 358456
rect 3846 358400 3851 358456
rect -960 358398 3851 358400
rect -960 358308 480 358398
rect 3785 358395 3851 358398
rect 238518 356628 238524 356692
rect 238588 356690 238594 356692
rect 238588 356630 240242 356690
rect 238588 356628 238594 356630
rect 240182 356080 240242 356630
rect 237373 355874 237439 355877
rect 237373 355872 240242 355874
rect 237373 355816 237378 355872
rect 237434 355816 240242 355872
rect 237373 355814 240242 355816
rect 237373 355811 237439 355814
rect 240182 355264 240242 355814
rect 237373 354650 237439 354653
rect 237373 354648 240242 354650
rect 237373 354592 237378 354648
rect 237434 354592 240242 354648
rect 237373 354590 240242 354592
rect 237373 354587 237439 354590
rect 240182 354312 240242 354590
rect 238334 351868 238340 351932
rect 238404 351930 238410 351932
rect 238404 351870 240242 351930
rect 238404 351868 238410 351870
rect 240182 351728 240242 351870
rect 583520 351780 584960 352020
rect 237373 351522 237439 351525
rect 237373 351520 240242 351522
rect 237373 351464 237378 351520
rect 237434 351464 240242 351520
rect 237373 351462 240242 351464
rect 237373 351459 237439 351462
rect 240182 350912 240242 351462
rect 237373 350298 237439 350301
rect 237373 350296 240242 350298
rect 237373 350240 237378 350296
rect 237434 350240 240242 350296
rect 237373 350238 240242 350240
rect 237373 350235 237439 350238
rect 240182 349960 240242 350238
rect 237373 347578 237439 347581
rect 237373 347576 240242 347578
rect 237373 347520 237378 347576
rect 237434 347520 240242 347576
rect 237373 347518 240242 347520
rect 237373 347515 237439 347518
rect 240182 347376 240242 347518
rect 237465 347034 237531 347037
rect 237465 347032 240242 347034
rect 237465 346976 237470 347032
rect 237526 346976 240242 347032
rect 237465 346974 240242 346976
rect 237465 346971 237531 346974
rect 240182 346424 240242 346974
rect 237373 346218 237439 346221
rect 237373 346216 240242 346218
rect 237373 346160 237378 346216
rect 237434 346160 240242 346216
rect 237373 346158 240242 346160
rect 237373 346155 237439 346158
rect 240182 345608 240242 346158
rect -960 345402 480 345492
rect -960 345342 6930 345402
rect -960 345252 480 345342
rect 6870 345130 6930 345342
rect 235206 345130 235212 345132
rect 6870 345070 235212 345130
rect 235206 345068 235212 345070
rect 235276 345068 235282 345132
rect 237373 343498 237439 343501
rect 237373 343496 240242 343498
rect 237373 343440 237378 343496
rect 237434 343440 240242 343496
rect 237373 343438 240242 343440
rect 237373 343435 237439 343438
rect 240182 343024 240242 343438
rect 237373 342138 237439 342141
rect 237373 342136 240242 342138
rect 237373 342080 237378 342136
rect 237434 342080 240242 342136
rect 237373 342078 240242 342080
rect 237373 342075 237439 342078
rect 240182 342072 240242 342078
rect 237465 341866 237531 341869
rect 237465 341864 240242 341866
rect 237465 341808 237470 341864
rect 237526 341808 240242 341864
rect 237465 341806 240242 341808
rect 237465 341803 237531 341806
rect 240182 341256 240242 341806
rect 237373 339146 237439 339149
rect 237373 339144 240242 339146
rect 237373 339088 237378 339144
rect 237434 339088 240242 339144
rect 237373 339086 240242 339088
rect 237373 339083 237439 339086
rect 240182 338536 240242 339086
rect 583520 338452 584960 338692
rect 237373 337922 237439 337925
rect 237373 337920 240242 337922
rect 237373 337864 237378 337920
rect 237434 337864 240242 337920
rect 237373 337862 240242 337864
rect 237373 337859 237439 337862
rect 240182 337720 240242 337862
rect 237465 337378 237531 337381
rect 237465 337376 240242 337378
rect 237465 337320 237470 337376
rect 237526 337320 240242 337376
rect 237465 337318 240242 337320
rect 237465 337315 237531 337318
rect 240182 336768 240242 337318
rect 237373 336562 237439 336565
rect 237373 336560 240242 336562
rect 237373 336504 237378 336560
rect 237434 336504 240242 336560
rect 237373 336502 240242 336504
rect 237373 336499 237439 336502
rect 240182 335952 240242 336502
rect 237373 335202 237439 335205
rect 237373 335200 240242 335202
rect 237373 335144 237378 335200
rect 237434 335144 240242 335200
rect 237373 335142 240242 335144
rect 237373 335139 237439 335142
rect 240182 335000 240242 335142
rect 237465 334794 237531 334797
rect 237465 334792 240242 334794
rect 237465 334736 237470 334792
rect 237526 334736 240242 334792
rect 237465 334734 240242 334736
rect 237465 334731 237531 334734
rect 240182 334184 240242 334734
rect 237373 333842 237439 333845
rect 237373 333840 240242 333842
rect 237373 333784 237378 333840
rect 237434 333784 240242 333840
rect 237373 333782 240242 333784
rect 237373 333779 237439 333782
rect 240182 333232 240242 333782
rect 237373 332482 237439 332485
rect 237373 332480 240242 332482
rect -960 332196 480 332436
rect 237373 332424 237378 332480
rect 237434 332424 240242 332480
rect 237373 332422 240242 332424
rect 237373 332419 237439 332422
rect 240182 332416 240242 332422
rect 237465 332210 237531 332213
rect 237465 332208 240242 332210
rect 237465 332152 237470 332208
rect 237526 332152 240242 332208
rect 237465 332150 240242 332152
rect 237465 332147 237531 332150
rect 240182 331600 240242 332150
rect 237373 330986 237439 330989
rect 237373 330984 240242 330986
rect 237373 330928 237378 330984
rect 237434 330928 240242 330984
rect 237373 330926 240242 330928
rect 237373 330923 237439 330926
rect 240182 330648 240242 330926
rect 238150 329700 238156 329764
rect 238220 329762 238226 329764
rect 240182 329762 240242 329776
rect 238220 329702 240242 329762
rect 238220 329700 238226 329702
rect 237373 329490 237439 329493
rect 237373 329488 240242 329490
rect 237373 329432 237378 329488
rect 237434 329432 240242 329488
rect 237373 329430 240242 329432
rect 237373 329427 237439 329430
rect 240182 328880 240242 329430
rect 237373 328266 237439 328269
rect 237373 328264 240242 328266
rect 237373 328208 237378 328264
rect 237434 328208 240242 328264
rect 237373 328206 240242 328208
rect 237373 328203 237439 328206
rect 240182 328064 240242 328206
rect 237465 327722 237531 327725
rect 237465 327720 240242 327722
rect 237465 327664 237470 327720
rect 237526 327664 240242 327720
rect 237465 327662 240242 327664
rect 237465 327659 237531 327662
rect 240182 327112 240242 327662
rect 237373 326906 237439 326909
rect 237373 326904 240242 326906
rect 237373 326848 237378 326904
rect 237434 326848 240242 326904
rect 237373 326846 240242 326848
rect 237373 326843 237439 326846
rect 240182 326296 240242 326846
rect 237465 325546 237531 325549
rect 237465 325544 240242 325546
rect 237465 325488 237470 325544
rect 237526 325488 240242 325544
rect 237465 325486 240242 325488
rect 237465 325483 237531 325486
rect 240182 325344 240242 325486
rect 579981 325274 580047 325277
rect 583520 325274 584960 325364
rect 579981 325272 584960 325274
rect 579981 325216 579986 325272
rect 580042 325216 584960 325272
rect 579981 325214 584960 325216
rect 579981 325211 580047 325214
rect 237373 325138 237439 325141
rect 237373 325136 240242 325138
rect 237373 325080 237378 325136
rect 237434 325080 240242 325136
rect 583520 325124 584960 325214
rect 237373 325078 240242 325080
rect 237373 325075 237439 325078
rect 240182 324528 240242 325078
rect 237373 324186 237439 324189
rect 237373 324184 240242 324186
rect 237373 324128 237378 324184
rect 237434 324128 240242 324184
rect 237373 324126 240242 324128
rect 237373 324123 237439 324126
rect 240182 323576 240242 324126
rect 237373 322826 237439 322829
rect 237373 322824 240242 322826
rect 237373 322768 237378 322824
rect 237434 322768 240242 322824
rect 237373 322766 240242 322768
rect 237373 322763 237439 322766
rect 240182 322760 240242 322766
rect 238293 322418 238359 322421
rect 238293 322416 240242 322418
rect 238293 322360 238298 322416
rect 238354 322360 240242 322416
rect 238293 322358 240242 322360
rect 238293 322355 238359 322358
rect 240182 321808 240242 322358
rect 237373 321466 237439 321469
rect 237373 321464 240242 321466
rect 237373 321408 237378 321464
rect 237434 321408 240242 321464
rect 237373 321406 240242 321408
rect 237373 321403 237439 321406
rect 240182 320992 240242 321406
rect 237373 320106 237439 320109
rect 240182 320106 240242 320120
rect 237373 320104 240242 320106
rect 237373 320048 237378 320104
rect 237434 320048 240242 320104
rect 237373 320046 240242 320048
rect 237373 320043 237439 320046
rect 237465 319834 237531 319837
rect 237465 319832 240242 319834
rect 237465 319776 237470 319832
rect 237526 319776 240242 319832
rect 237465 319774 240242 319776
rect 237465 319771 237531 319774
rect -960 319140 480 319380
rect 240182 319224 240242 319774
rect 237373 318610 237439 318613
rect 237373 318608 240242 318610
rect 237373 318552 237378 318608
rect 237434 318552 240242 318608
rect 237373 318550 240242 318552
rect 237373 318547 237439 318550
rect 240182 318408 240242 318550
rect 238017 318066 238083 318069
rect 238017 318064 240242 318066
rect 238017 318008 238022 318064
rect 238078 318008 240242 318064
rect 238017 318006 240242 318008
rect 238017 318003 238083 318006
rect 240182 317456 240242 318006
rect 237373 317250 237439 317253
rect 237373 317248 240242 317250
rect 237373 317192 237378 317248
rect 237434 317192 240242 317248
rect 237373 317190 240242 317192
rect 237373 317187 237439 317190
rect 240182 316640 240242 317190
rect 237966 315964 237972 316028
rect 238036 316026 238042 316028
rect 238036 315966 240242 316026
rect 238036 315964 238042 315966
rect 240182 315688 240242 315966
rect 237373 315482 237439 315485
rect 237373 315480 240242 315482
rect 237373 315424 237378 315480
rect 237434 315424 240242 315480
rect 237373 315422 240242 315424
rect 237373 315419 237439 315422
rect 240182 314872 240242 315422
rect 237373 314530 237439 314533
rect 237373 314528 240242 314530
rect 237373 314472 237378 314528
rect 237434 314472 240242 314528
rect 237373 314470 240242 314472
rect 237373 314467 237439 314470
rect 240182 313920 240242 314470
rect 237373 313170 237439 313173
rect 237373 313168 240242 313170
rect 237373 313112 237378 313168
rect 237434 313112 240242 313168
rect 237373 313110 240242 313112
rect 237373 313107 237439 313110
rect 240182 313104 240242 313110
rect 237465 312762 237531 312765
rect 237465 312760 240242 312762
rect 237465 312704 237470 312760
rect 237526 312704 240242 312760
rect 237465 312702 240242 312704
rect 237465 312699 237531 312702
rect 240182 312152 240242 312702
rect 580165 312082 580231 312085
rect 583520 312082 584960 312172
rect 580165 312080 584960 312082
rect 580165 312024 580170 312080
rect 580226 312024 584960 312080
rect 580165 312022 584960 312024
rect 580165 312019 580231 312022
rect 583520 311932 584960 312022
rect 237373 311810 237439 311813
rect 237373 311808 240242 311810
rect 237373 311752 237378 311808
rect 237434 311752 240242 311808
rect 237373 311750 240242 311752
rect 237373 311747 237439 311750
rect 240182 311336 240242 311750
rect 237373 310450 237439 310453
rect 240182 310450 240242 310464
rect 237373 310448 240242 310450
rect 237373 310392 237378 310448
rect 237434 310392 240242 310448
rect 237373 310390 240242 310392
rect 237373 310387 237439 310390
rect 237465 310178 237531 310181
rect 237465 310176 240242 310178
rect 237465 310120 237470 310176
rect 237526 310120 240242 310176
rect 237465 310118 240242 310120
rect 237465 310115 237531 310118
rect 240182 309568 240242 310118
rect 237373 308954 237439 308957
rect 237373 308952 240242 308954
rect 237373 308896 237378 308952
rect 237434 308896 240242 308952
rect 237373 308894 240242 308896
rect 237373 308891 237439 308894
rect 240182 308752 240242 308894
rect 237465 308410 237531 308413
rect 237465 308408 240242 308410
rect 237465 308352 237470 308408
rect 237526 308352 240242 308408
rect 237465 308350 240242 308352
rect 237465 308347 237531 308350
rect 240182 307800 240242 308350
rect 237373 307594 237439 307597
rect 237373 307592 240242 307594
rect 237373 307536 237378 307592
rect 237434 307536 240242 307592
rect 237373 307534 240242 307536
rect 237373 307531 237439 307534
rect 240182 306984 240242 307534
rect -960 306234 480 306324
rect 3141 306234 3207 306237
rect -960 306232 3207 306234
rect -960 306176 3146 306232
rect 3202 306176 3207 306232
rect -960 306174 3207 306176
rect -960 306084 480 306174
rect 3141 306171 3207 306174
rect 237373 306234 237439 306237
rect 237373 306232 240242 306234
rect 237373 306176 237378 306232
rect 237434 306176 240242 306232
rect 237373 306174 240242 306176
rect 237373 306171 237439 306174
rect 240182 306032 240242 306174
rect 237465 305826 237531 305829
rect 237465 305824 240242 305826
rect 237465 305768 237470 305824
rect 237526 305768 240242 305824
rect 237465 305766 240242 305768
rect 237465 305763 237531 305766
rect 240182 305216 240242 305766
rect 237373 304874 237439 304877
rect 237373 304872 240242 304874
rect 237373 304816 237378 304872
rect 237434 304816 240242 304872
rect 237373 304814 240242 304816
rect 237373 304811 237439 304814
rect 240182 304264 240242 304814
rect 237373 303514 237439 303517
rect 237373 303512 240242 303514
rect 237373 303456 237378 303512
rect 237434 303456 240242 303512
rect 237373 303454 240242 303456
rect 237373 303451 237439 303454
rect 240182 303448 240242 303454
rect 237465 303106 237531 303109
rect 237465 303104 240242 303106
rect 237465 303048 237470 303104
rect 237526 303048 240242 303104
rect 237465 303046 240242 303048
rect 237465 303043 237531 303046
rect 240182 302496 240242 303046
rect 237373 302154 237439 302157
rect 237373 302152 240242 302154
rect 237373 302096 237378 302152
rect 237434 302096 240242 302152
rect 237373 302094 240242 302096
rect 237373 302091 237439 302094
rect 240182 301680 240242 302094
rect 237373 300794 237439 300797
rect 237373 300792 240242 300794
rect 237373 300736 237378 300792
rect 237434 300736 240242 300792
rect 237373 300734 240242 300736
rect 237373 300731 237439 300734
rect 240182 300728 240242 300734
rect 237465 300522 237531 300525
rect 237465 300520 240242 300522
rect 237465 300464 237470 300520
rect 237526 300464 240242 300520
rect 237465 300462 240242 300464
rect 237465 300459 237531 300462
rect 240182 299912 240242 300462
rect 237373 299298 237439 299301
rect 237373 299296 240242 299298
rect 237373 299240 237378 299296
rect 237434 299240 240242 299296
rect 237373 299238 240242 299240
rect 237373 299235 237439 299238
rect 240182 299096 240242 299238
rect 237465 298754 237531 298757
rect 237465 298752 240242 298754
rect 237465 298696 237470 298752
rect 237526 298696 240242 298752
rect 237465 298694 240242 298696
rect 237465 298691 237531 298694
rect 240182 298144 240242 298694
rect 583520 298604 584960 298844
rect 237373 297938 237439 297941
rect 237373 297936 240242 297938
rect 237373 297880 237378 297936
rect 237434 297880 240242 297936
rect 237373 297878 240242 297880
rect 237373 297875 237439 297878
rect 240182 297328 240242 297878
rect 237373 296578 237439 296581
rect 237373 296576 240242 296578
rect 237373 296520 237378 296576
rect 237434 296520 240242 296576
rect 237373 296518 240242 296520
rect 237373 296515 237439 296518
rect 240182 296376 240242 296518
rect 237465 296170 237531 296173
rect 237465 296168 240242 296170
rect 237465 296112 237470 296168
rect 237526 296112 240242 296168
rect 237465 296110 240242 296112
rect 237465 296107 237531 296110
rect 240182 295560 240242 296110
rect 237373 295218 237439 295221
rect 237373 295216 240242 295218
rect 237373 295160 237378 295216
rect 237434 295160 240242 295216
rect 237373 295158 240242 295160
rect 237373 295155 237439 295158
rect 240182 294608 240242 295158
rect 237373 293858 237439 293861
rect 237373 293856 240242 293858
rect 237373 293800 237378 293856
rect 237434 293800 240242 293856
rect 237373 293798 240242 293800
rect 237373 293795 237439 293798
rect 240182 293792 240242 293798
rect -960 293178 480 293268
rect 3325 293178 3391 293181
rect -960 293176 3391 293178
rect -960 293120 3330 293176
rect 3386 293120 3391 293176
rect -960 293118 3391 293120
rect -960 293028 480 293118
rect 3325 293115 3391 293118
rect 237373 292770 237439 292773
rect 240182 292770 240242 292784
rect 237373 292768 240242 292770
rect 237373 292712 237378 292768
rect 237434 292712 240242 292768
rect 237373 292710 240242 292712
rect 237373 292707 237439 292710
rect 237373 291410 237439 291413
rect 240182 291410 240242 291968
rect 237373 291408 240242 291410
rect 237373 291352 237378 291408
rect 237434 291352 240242 291408
rect 237373 291350 240242 291352
rect 237373 291347 237439 291350
rect 235574 290396 235580 290460
rect 235644 290458 235650 290460
rect 240182 290458 240242 291016
rect 235644 290398 240242 290458
rect 235644 290396 235650 290398
rect 237373 290050 237439 290053
rect 240182 290050 240242 290200
rect 237373 290048 240242 290050
rect 237373 289992 237378 290048
rect 237434 289992 240242 290048
rect 237373 289990 240242 289992
rect 237373 289987 237439 289990
rect 237465 288690 237531 288693
rect 240182 288690 240242 289248
rect 237465 288688 240242 288690
rect 237465 288632 237470 288688
rect 237526 288632 240242 288688
rect 237465 288630 240242 288632
rect 237465 288627 237531 288630
rect 237373 288554 237439 288557
rect 237373 288552 240242 288554
rect 237373 288496 237378 288552
rect 237434 288496 240242 288552
rect 237373 288494 240242 288496
rect 237373 288491 237439 288494
rect 240182 288488 240242 288494
rect 237373 287194 237439 287197
rect 240182 287194 240242 287616
rect 237373 287192 240242 287194
rect 237373 287136 237378 287192
rect 237434 287136 240242 287192
rect 237373 287134 240242 287136
rect 237373 287131 237439 287134
rect 49601 286378 49667 286381
rect 180701 286378 180767 286381
rect 49601 286376 180767 286378
rect 49601 286320 49606 286376
rect 49662 286320 180706 286376
rect 180762 286320 180767 286376
rect 49601 286318 180767 286320
rect 49601 286315 49667 286318
rect 180701 286315 180767 286318
rect 136030 286180 136036 286244
rect 136100 286242 136106 286244
rect 136541 286242 136607 286245
rect 136100 286240 136607 286242
rect 136100 286184 136546 286240
rect 136602 286184 136607 286240
rect 136100 286182 136607 286184
rect 136100 286180 136106 286182
rect 136541 286179 136607 286182
rect 138422 286180 138428 286244
rect 138492 286242 138498 286244
rect 139301 286242 139367 286245
rect 138492 286240 139367 286242
rect 138492 286184 139306 286240
rect 139362 286184 139367 286240
rect 138492 286182 139367 286184
rect 138492 286180 138498 286182
rect 139301 286179 139367 286182
rect 143574 286180 143580 286244
rect 143644 286242 143650 286244
rect 144821 286242 144887 286245
rect 143644 286240 144887 286242
rect 143644 286184 144826 286240
rect 144882 286184 144887 286240
rect 143644 286182 144887 286184
rect 143644 286180 143650 286182
rect 144821 286179 144887 286182
rect 169702 286180 169708 286244
rect 169772 286242 169778 286244
rect 170673 286242 170739 286245
rect 169772 286240 170739 286242
rect 169772 286184 170678 286240
rect 170734 286184 170739 286240
rect 169772 286182 170739 286184
rect 169772 286180 169778 286182
rect 170673 286179 170739 286182
rect 78806 286044 78812 286108
rect 78876 286106 78882 286108
rect 235390 286106 235396 286108
rect 78876 286046 235396 286106
rect 78876 286044 78882 286046
rect 235390 286044 235396 286046
rect 235460 286044 235466 286108
rect 237373 286106 237439 286109
rect 240182 286106 240242 286664
rect 237373 286104 240242 286106
rect 237373 286048 237378 286104
rect 237434 286048 240242 286104
rect 237373 286046 240242 286048
rect 237373 286043 237439 286046
rect 106181 285972 106247 285973
rect 106181 285970 106228 285972
rect 106136 285968 106228 285970
rect 106136 285912 106186 285968
rect 106136 285910 106228 285912
rect 106181 285908 106228 285910
rect 106292 285908 106298 285972
rect 108430 285908 108436 285972
rect 108500 285970 108506 285972
rect 108941 285970 109007 285973
rect 108500 285968 109007 285970
rect 108500 285912 108946 285968
rect 109002 285912 109007 285968
rect 108500 285910 109007 285912
rect 108500 285908 108506 285910
rect 106181 285907 106247 285908
rect 108941 285907 109007 285910
rect 120758 285908 120764 285972
rect 120828 285970 120834 285972
rect 187182 285970 187188 285972
rect 120828 285910 187188 285970
rect 120828 285908 120834 285910
rect 187182 285908 187188 285910
rect 187252 285908 187258 285972
rect 81014 285772 81020 285836
rect 81084 285834 81090 285836
rect 232497 285834 232563 285837
rect 81084 285832 232563 285834
rect 81084 285776 232502 285832
rect 232558 285776 232563 285832
rect 81084 285774 232563 285776
rect 81084 285772 81090 285774
rect 232497 285771 232563 285774
rect 237465 285834 237531 285837
rect 240182 285834 240242 285848
rect 237465 285832 240242 285834
rect 237465 285776 237470 285832
rect 237526 285776 240242 285832
rect 237465 285774 240242 285776
rect 237465 285771 237531 285774
rect 83406 285636 83412 285700
rect 83476 285698 83482 285700
rect 83733 285698 83799 285701
rect 83476 285696 83799 285698
rect 83476 285640 83738 285696
rect 83794 285640 83799 285696
rect 83476 285638 83799 285640
rect 83476 285636 83482 285638
rect 83733 285635 83799 285638
rect 86166 285636 86172 285700
rect 86236 285698 86242 285700
rect 86861 285698 86927 285701
rect 86236 285696 86927 285698
rect 86236 285640 86866 285696
rect 86922 285640 86927 285696
rect 86236 285638 86927 285640
rect 86236 285636 86242 285638
rect 86861 285635 86927 285638
rect 88558 285636 88564 285700
rect 88628 285698 88634 285700
rect 89621 285698 89687 285701
rect 88628 285696 89687 285698
rect 88628 285640 89626 285696
rect 89682 285640 89687 285696
rect 88628 285638 89687 285640
rect 88628 285636 88634 285638
rect 89621 285635 89687 285638
rect 91134 285636 91140 285700
rect 91204 285698 91210 285700
rect 92381 285698 92447 285701
rect 91204 285696 92447 285698
rect 91204 285640 92386 285696
rect 92442 285640 92447 285696
rect 91204 285638 92447 285640
rect 91204 285636 91210 285638
rect 92381 285635 92447 285638
rect 93526 285636 93532 285700
rect 93596 285698 93602 285700
rect 93669 285698 93735 285701
rect 93596 285696 93735 285698
rect 93596 285640 93674 285696
rect 93730 285640 93735 285696
rect 93596 285638 93735 285640
rect 93596 285636 93602 285638
rect 93669 285635 93735 285638
rect 96286 285636 96292 285700
rect 96356 285698 96362 285700
rect 96521 285698 96587 285701
rect 96356 285696 96587 285698
rect 96356 285640 96526 285696
rect 96582 285640 96587 285696
rect 96356 285638 96587 285640
rect 96356 285636 96362 285638
rect 96521 285635 96587 285638
rect 103830 285636 103836 285700
rect 103900 285698 103906 285700
rect 104801 285698 104867 285701
rect 103900 285696 104867 285698
rect 103900 285640 104806 285696
rect 104862 285640 104867 285696
rect 103900 285638 104867 285640
rect 103900 285636 103906 285638
rect 104801 285635 104867 285638
rect 114318 285636 114324 285700
rect 114388 285698 114394 285700
rect 114461 285698 114527 285701
rect 118601 285700 118667 285701
rect 114388 285696 114527 285698
rect 114388 285640 114466 285696
rect 114522 285640 114527 285696
rect 114388 285638 114527 285640
rect 114388 285636 114394 285638
rect 114461 285635 114527 285638
rect 118550 285636 118556 285700
rect 118620 285698 118667 285700
rect 118620 285696 118712 285698
rect 118662 285640 118712 285696
rect 118620 285638 118712 285640
rect 118620 285636 118667 285638
rect 123518 285636 123524 285700
rect 123588 285698 123594 285700
rect 124121 285698 124187 285701
rect 123588 285696 124187 285698
rect 123588 285640 124126 285696
rect 124182 285640 124187 285696
rect 123588 285638 124187 285640
rect 123588 285636 123594 285638
rect 118601 285635 118667 285636
rect 124121 285635 124187 285638
rect 125910 285636 125916 285700
rect 125980 285698 125986 285700
rect 126881 285698 126947 285701
rect 125980 285696 126947 285698
rect 125980 285640 126886 285696
rect 126942 285640 126947 285696
rect 125980 285638 126947 285640
rect 125980 285636 125986 285638
rect 126881 285635 126947 285638
rect 133454 285636 133460 285700
rect 133524 285698 133530 285700
rect 133781 285698 133847 285701
rect 133524 285696 133847 285698
rect 133524 285640 133786 285696
rect 133842 285640 133847 285696
rect 133524 285638 133847 285640
rect 133524 285636 133530 285638
rect 133781 285635 133847 285638
rect 140998 285636 141004 285700
rect 141068 285698 141074 285700
rect 141877 285698 141943 285701
rect 141068 285696 141943 285698
rect 141068 285640 141882 285696
rect 141938 285640 141943 285696
rect 141068 285638 141943 285640
rect 141068 285636 141074 285638
rect 141877 285635 141943 285638
rect 151118 285636 151124 285700
rect 151188 285698 151194 285700
rect 151721 285698 151787 285701
rect 151188 285696 151787 285698
rect 151188 285640 151726 285696
rect 151782 285640 151787 285696
rect 151188 285638 151787 285640
rect 151188 285636 151194 285638
rect 151721 285635 151787 285638
rect 154062 285636 154068 285700
rect 154132 285698 154138 285700
rect 154481 285698 154547 285701
rect 154132 285696 154547 285698
rect 154132 285640 154486 285696
rect 154542 285640 154547 285696
rect 154132 285638 154547 285640
rect 154132 285636 154138 285638
rect 154481 285635 154547 285638
rect 156086 285636 156092 285700
rect 156156 285698 156162 285700
rect 157241 285698 157307 285701
rect 156156 285696 157307 285698
rect 156156 285640 157246 285696
rect 157302 285640 157307 285696
rect 156156 285638 157307 285640
rect 156156 285636 156162 285638
rect 157241 285635 157307 285638
rect 168414 285636 168420 285700
rect 168484 285698 168490 285700
rect 169661 285698 169727 285701
rect 168484 285696 169727 285698
rect 168484 285640 169666 285696
rect 169722 285640 169727 285696
rect 168484 285638 169727 285640
rect 168484 285636 168490 285638
rect 169661 285635 169727 285638
rect 583520 285276 584960 285516
rect 128721 285156 128787 285157
rect 131113 285156 131179 285157
rect 128670 285092 128676 285156
rect 128740 285154 128787 285156
rect 128740 285152 128832 285154
rect 128782 285096 128832 285152
rect 128740 285094 128832 285096
rect 128740 285092 128787 285094
rect 131062 285092 131068 285156
rect 131132 285154 131179 285156
rect 131132 285152 131224 285154
rect 131174 285096 131224 285152
rect 131132 285094 131224 285096
rect 131132 285092 131179 285094
rect 128721 285091 128787 285092
rect 131113 285091 131179 285092
rect 111057 285020 111123 285021
rect 116209 285020 116275 285021
rect 111006 284956 111012 285020
rect 111076 285018 111123 285020
rect 111076 285016 111168 285018
rect 111118 284960 111168 285016
rect 111076 284958 111168 284960
rect 111076 284956 111123 284958
rect 116158 284956 116164 285020
rect 116228 285018 116275 285020
rect 116228 285016 116320 285018
rect 116270 284960 116320 285016
rect 116228 284958 116320 284960
rect 116228 284956 116275 284958
rect 111057 284955 111123 284956
rect 116209 284955 116275 284956
rect 98545 284884 98611 284885
rect 148593 284884 148659 284885
rect 98494 284820 98500 284884
rect 98564 284882 98611 284884
rect 98564 284880 98656 284882
rect 98606 284824 98656 284880
rect 98564 284822 98656 284824
rect 98564 284820 98611 284822
rect 148542 284820 148548 284884
rect 148612 284882 148659 284884
rect 237373 284882 237439 284885
rect 240182 284882 240242 284896
rect 148612 284880 148704 284882
rect 148654 284824 148704 284880
rect 148612 284822 148704 284824
rect 237373 284880 240242 284882
rect 237373 284824 237378 284880
rect 237434 284824 240242 284880
rect 237373 284822 240242 284824
rect 148612 284820 148659 284822
rect 98545 284819 98611 284820
rect 148593 284819 148659 284820
rect 237373 284819 237439 284822
rect 101305 284748 101371 284749
rect 146017 284748 146083 284749
rect 101254 284684 101260 284748
rect 101324 284746 101371 284748
rect 101324 284744 101416 284746
rect 101366 284688 101416 284744
rect 101324 284686 101416 284688
rect 101324 284684 101371 284686
rect 145966 284684 145972 284748
rect 146036 284746 146083 284748
rect 146036 284744 146128 284746
rect 146078 284688 146128 284744
rect 146036 284686 146128 284688
rect 146036 284684 146083 284686
rect 101305 284683 101371 284684
rect 146017 284683 146083 284684
rect 180701 284068 180767 284069
rect 180701 284066 180748 284068
rect 180656 284064 180748 284066
rect 180812 284066 180818 284068
rect 180656 284008 180706 284064
rect 180656 284006 180748 284008
rect 180701 284004 180748 284006
rect 180812 284006 180894 284066
rect 180812 284004 180818 284006
rect 180701 284003 180767 284004
rect 237373 283522 237439 283525
rect 240182 283522 240242 284080
rect 237373 283520 240242 283522
rect 237373 283464 237378 283520
rect 237434 283464 240242 283520
rect 237373 283462 240242 283464
rect 237373 283459 237439 283462
rect 237465 282978 237531 282981
rect 240182 282978 240242 283128
rect 237465 282976 240242 282978
rect 237465 282920 237470 282976
rect 237526 282920 240242 282976
rect 237465 282918 240242 282920
rect 237465 282915 237531 282918
rect 237373 282842 237439 282845
rect 237373 282840 240242 282842
rect 237373 282784 237378 282840
rect 237434 282784 240242 282840
rect 237373 282782 240242 282784
rect 237373 282779 237439 282782
rect 240182 282368 240242 282782
rect 237373 280802 237439 280805
rect 240182 280802 240242 281360
rect 237373 280800 240242 280802
rect 237373 280744 237378 280800
rect 237434 280744 240242 280800
rect 237373 280742 240242 280744
rect 237373 280739 237439 280742
rect 237465 280394 237531 280397
rect 240182 280394 240242 280544
rect 237465 280392 240242 280394
rect 237465 280336 237470 280392
rect 237526 280336 240242 280392
rect 237465 280334 240242 280336
rect 237465 280331 237531 280334
rect -960 279972 480 280212
rect 237373 279850 237439 279853
rect 237373 279848 240242 279850
rect 237373 279792 237378 279848
rect 237434 279792 240242 279848
rect 237373 279790 240242 279792
rect 237373 279787 237439 279790
rect 240182 279648 240242 279790
rect 186588 279170 187250 279220
rect 189993 279170 190059 279173
rect 186588 279168 190059 279170
rect 186588 279160 189998 279168
rect 187190 279112 189998 279160
rect 190054 279112 190059 279168
rect 187190 279110 190059 279112
rect 189993 279107 190059 279110
rect 188286 278972 188292 279036
rect 188356 279034 188362 279036
rect 188356 278974 240242 279034
rect 188356 278972 188362 278974
rect 240182 278832 240242 278974
rect 186814 277476 186820 277540
rect 186884 277538 186890 277540
rect 240182 277538 240242 277960
rect 186884 277478 240242 277538
rect 186884 277476 186890 277478
rect 237373 277266 237439 277269
rect 237373 277264 240242 277266
rect 237373 277208 237378 277264
rect 237434 277208 240242 277264
rect 237373 277206 240242 277208
rect 237373 277203 237439 277206
rect 240182 277064 240242 277206
rect 188470 276116 188476 276180
rect 188540 276178 188546 276180
rect 240182 276178 240242 276192
rect 188540 276118 240242 276178
rect 188540 276116 188546 276118
rect 237465 275090 237531 275093
rect 240182 275090 240242 275240
rect 237465 275088 240242 275090
rect 237465 275032 237470 275088
rect 237526 275032 240242 275088
rect 237465 275030 240242 275032
rect 237465 275027 237531 275030
rect 237373 274546 237439 274549
rect 237373 274544 240242 274546
rect 237373 274488 237378 274544
rect 237434 274488 240242 274544
rect 237373 274486 240242 274488
rect 237373 274483 237439 274486
rect 240182 274480 240242 274486
rect 188654 273396 188660 273460
rect 188724 273458 188730 273460
rect 240182 273458 240242 273472
rect 188724 273398 240242 273458
rect 188724 273396 188730 273398
rect 186998 271900 187004 271964
rect 187068 271962 187074 271964
rect 240182 271962 240242 272656
rect 579797 272234 579863 272237
rect 583520 272234 584960 272324
rect 579797 272232 584960 272234
rect 579797 272176 579802 272232
rect 579858 272176 584960 272232
rect 579797 272174 584960 272176
rect 579797 272171 579863 272174
rect 583520 272084 584960 272174
rect 187068 271902 240242 271962
rect 187068 271900 187074 271902
rect 237373 271826 237439 271829
rect 237373 271824 240242 271826
rect 237373 271768 237378 271824
rect 237434 271768 240242 271824
rect 237373 271766 240242 271768
rect 237373 271763 237439 271766
rect 240182 271760 240242 271766
rect 238293 270738 238359 270741
rect 240182 270738 240242 270888
rect 238293 270736 240242 270738
rect 238293 270680 238298 270736
rect 238354 270680 240242 270736
rect 238293 270678 240242 270680
rect 238293 270675 238359 270678
rect 237966 269860 237972 269924
rect 238036 269922 238042 269924
rect 240182 269922 240242 269936
rect 238036 269862 240242 269922
rect 238036 269860 238042 269862
rect 237833 269786 237899 269789
rect 237833 269784 240242 269786
rect 237833 269728 237838 269784
rect 237894 269728 240242 269784
rect 237833 269726 240242 269728
rect 237833 269723 237899 269726
rect 240182 269176 240242 269726
rect 237373 267882 237439 267885
rect 240182 267882 240242 268168
rect 237373 267880 240242 267882
rect 237373 267824 237378 267880
rect 237434 267824 240242 267880
rect 237373 267822 240242 267824
rect 237373 267819 237439 267822
rect -960 267052 480 267292
rect 238150 267276 238156 267340
rect 238220 267338 238226 267340
rect 240182 267338 240242 267352
rect 238220 267278 240242 267338
rect 238220 267276 238226 267278
rect 238477 267202 238543 267205
rect 238477 267200 240242 267202
rect 238477 267144 238482 267200
rect 238538 267144 240242 267200
rect 238477 267142 240242 267144
rect 238477 267139 238543 267142
rect 240182 266592 240242 267142
rect 238477 265026 238543 265029
rect 240182 265026 240242 265584
rect 238477 265024 240242 265026
rect 238477 264968 238482 265024
rect 238538 264968 240242 265024
rect 238477 264966 240242 264968
rect 238477 264963 238543 264966
rect 238334 264148 238340 264212
rect 238404 264210 238410 264212
rect 240182 264210 240242 264768
rect 238404 264150 240242 264210
rect 238404 264148 238410 264150
rect 238661 264074 238727 264077
rect 238661 264072 240242 264074
rect 238661 264016 238666 264072
rect 238722 264016 240242 264072
rect 238661 264014 240242 264016
rect 238661 264011 238727 264014
rect 240182 263872 240242 264014
rect 237373 262442 237439 262445
rect 240182 262442 240242 263000
rect 237373 262440 240242 262442
rect 237373 262384 237378 262440
rect 237434 262384 240242 262440
rect 237373 262382 240242 262384
rect 237373 262379 237439 262382
rect 237373 262034 237439 262037
rect 240182 262034 240242 262048
rect 237373 262032 240242 262034
rect 237373 261976 237378 262032
rect 237434 261976 240242 262032
rect 237373 261974 240242 261976
rect 237373 261971 237439 261974
rect 237465 261898 237531 261901
rect 237465 261896 240242 261898
rect 237465 261840 237470 261896
rect 237526 261840 240242 261896
rect 237465 261838 240242 261840
rect 237465 261835 237531 261838
rect 240182 261288 240242 261838
rect 237373 259722 237439 259725
rect 240182 259722 240242 260280
rect 237373 259720 240242 259722
rect 237373 259664 237378 259720
rect 237434 259664 240242 259720
rect 237373 259662 240242 259664
rect 237373 259659 237439 259662
rect 237465 259586 237531 259589
rect 237465 259584 240242 259586
rect 237465 259528 237470 259584
rect 237526 259528 240242 259584
rect 237465 259526 240242 259528
rect 237465 259523 237531 259526
rect 240182 259520 240242 259526
rect 237373 259178 237439 259181
rect 237373 259176 240242 259178
rect 237373 259120 237378 259176
rect 237434 259120 240242 259176
rect 237373 259118 240242 259120
rect 237373 259115 237439 259118
rect 240182 258568 240242 259118
rect 579981 258906 580047 258909
rect 583520 258906 584960 258996
rect 579981 258904 584960 258906
rect 579981 258848 579986 258904
rect 580042 258848 584960 258904
rect 579981 258846 584960 258848
rect 579981 258843 580047 258846
rect 583520 258756 584960 258846
rect 237373 257138 237439 257141
rect 240182 257138 240242 257696
rect 237373 257136 240242 257138
rect 237373 257080 237378 257136
rect 237434 257080 240242 257136
rect 237373 257078 240242 257080
rect 237373 257075 237439 257078
rect 237465 256866 237531 256869
rect 237465 256864 240242 256866
rect 237465 256808 237470 256864
rect 237526 256808 240242 256864
rect 237465 256806 240242 256808
rect 237465 256803 237531 256806
rect 240182 256800 240242 256806
rect 187182 255308 187188 255372
rect 187252 255370 187258 255372
rect 240182 255370 240242 255928
rect 187252 255310 240242 255370
rect 187252 255308 187258 255310
rect 237465 254554 237531 254557
rect 240182 254554 240242 255112
rect 237465 254552 240242 254554
rect 237465 254496 237470 254552
rect 237526 254496 240242 254552
rect 237465 254494 240242 254496
rect 237465 254491 237531 254494
rect -960 254146 480 254236
rect 2773 254146 2839 254149
rect -960 254144 2839 254146
rect -960 254088 2778 254144
rect 2834 254088 2839 254144
rect -960 254086 2839 254088
rect -960 253996 480 254086
rect 2773 254083 2839 254086
rect 237373 254146 237439 254149
rect 240182 254146 240242 254160
rect 237373 254144 240242 254146
rect 237373 254088 237378 254144
rect 237434 254088 240242 254144
rect 237373 254086 240242 254088
rect 237373 254083 237439 254086
rect 238109 253874 238175 253877
rect 238109 253872 240242 253874
rect 238109 253816 238114 253872
rect 238170 253816 240242 253872
rect 238109 253814 240242 253816
rect 238109 253811 238175 253814
rect 240182 253400 240242 253814
rect 237373 251834 237439 251837
rect 240182 251834 240242 252392
rect 237373 251832 240242 251834
rect 237373 251776 237378 251832
rect 237434 251776 240242 251832
rect 237373 251774 240242 251776
rect 237373 251771 237439 251774
rect 238109 251426 238175 251429
rect 240182 251426 240242 251576
rect 238109 251424 240242 251426
rect 238109 251368 238114 251424
rect 238170 251368 240242 251424
rect 238109 251366 240242 251368
rect 238109 251363 238175 251366
rect 238569 250882 238635 250885
rect 238569 250880 240242 250882
rect 238569 250824 238574 250880
rect 238630 250824 240242 250880
rect 238569 250822 240242 250824
rect 238569 250819 238635 250822
rect 240182 250680 240242 250822
rect 237373 249930 237439 249933
rect 237373 249928 240242 249930
rect 237373 249872 237378 249928
rect 237434 249872 240242 249928
rect 237373 249870 240242 249872
rect 237373 249867 237439 249870
rect 240182 249864 240242 249870
rect 237373 248570 237439 248573
rect 240182 248570 240242 248856
rect 237373 248568 240242 248570
rect 237373 248512 237378 248568
rect 237434 248512 240242 248568
rect 237373 248510 240242 248512
rect 237373 248507 237439 248510
rect 238201 248298 238267 248301
rect 238201 248296 240242 248298
rect 238201 248240 238206 248296
rect 238262 248240 240242 248296
rect 238201 248238 240242 248240
rect 238201 248235 238267 248238
rect 240182 248096 240242 248238
rect 237373 247074 237439 247077
rect 240182 247074 240242 247088
rect 237373 247072 240242 247074
rect 237373 247016 237378 247072
rect 237434 247016 240242 247072
rect 237373 247014 240242 247016
rect 237373 247011 237439 247014
rect 238201 245714 238267 245717
rect 240182 245714 240242 246272
rect 238201 245712 240242 245714
rect 238201 245656 238206 245712
rect 238262 245656 240242 245712
rect 238201 245654 240242 245656
rect 238201 245651 238267 245654
rect 238385 245578 238451 245581
rect 238385 245576 240242 245578
rect 238385 245520 238390 245576
rect 238446 245520 240242 245576
rect 238385 245518 240242 245520
rect 238385 245515 238451 245518
rect 240182 245512 240242 245518
rect 583520 245428 584960 245668
rect 237373 244490 237439 244493
rect 240182 244490 240242 244504
rect 237373 244488 240242 244490
rect 237373 244432 237378 244488
rect 237434 244432 240242 244488
rect 237373 244430 240242 244432
rect 237373 244427 237439 244430
rect 238385 243130 238451 243133
rect 240182 243130 240242 243688
rect 238385 243128 240242 243130
rect 238385 243072 238390 243128
rect 238446 243072 240242 243128
rect 238385 243070 240242 243072
rect 238385 243067 238451 243070
rect 237373 242858 237439 242861
rect 237373 242856 240242 242858
rect 237373 242800 237378 242856
rect 237434 242800 240242 242856
rect 237373 242798 240242 242800
rect 237373 242795 237439 242798
rect 240182 242792 240242 242798
rect 237373 241634 237439 241637
rect 240182 241634 240242 241920
rect 237373 241632 240242 241634
rect 237373 241576 237378 241632
rect 237434 241576 240242 241632
rect 237373 241574 240242 241576
rect 237373 241571 237439 241574
rect -960 241090 480 241180
rect 3141 241090 3207 241093
rect -960 241088 3207 241090
rect -960 241032 3146 241088
rect 3202 241032 3207 241088
rect -960 241030 3207 241032
rect -960 240940 480 241030
rect 3141 241027 3207 241030
rect 237373 240410 237439 240413
rect 240182 240410 240242 240968
rect 237373 240408 240242 240410
rect 237373 240352 237378 240408
rect 237434 240352 240242 240408
rect 237373 240350 240242 240352
rect 237373 240347 237439 240350
rect 237373 238642 237439 238645
rect 237373 238640 240242 238642
rect 237373 238584 237378 238640
rect 237434 238584 240242 238640
rect 237373 238582 240242 238584
rect 237373 238579 237439 238582
rect 240182 238440 240242 238582
rect 238569 237418 238635 237421
rect 240182 237418 240242 237432
rect 238569 237416 240242 237418
rect 238569 237360 238574 237416
rect 238630 237360 240242 237416
rect 238569 237358 240242 237360
rect 238569 237355 238635 237358
rect 48129 236874 48195 236877
rect 49374 236874 50048 236924
rect 48129 236872 50048 236874
rect 48129 236816 48134 236872
rect 48190 236864 50048 236872
rect 48190 236816 49434 236864
rect 48129 236814 49434 236816
rect 48129 236811 48195 236814
rect 237373 236058 237439 236061
rect 240182 236058 240242 236616
rect 237373 236056 240242 236058
rect 237373 236000 237378 236056
rect 237434 236000 240242 236056
rect 237373 235998 240242 236000
rect 237373 235995 237439 235998
rect 47945 235922 48011 235925
rect 49374 235922 50048 235972
rect 47945 235920 50048 235922
rect 47945 235864 47950 235920
rect 48006 235912 50048 235920
rect 48006 235864 49434 235912
rect 47945 235862 49434 235864
rect 47945 235859 48011 235862
rect 237373 234290 237439 234293
rect 237373 234288 240242 234290
rect 237373 234232 237378 234288
rect 237434 234232 240242 234288
rect 237373 234230 240242 234232
rect 237373 234227 237439 234230
rect 240182 234088 240242 234230
rect 47853 233746 47919 233749
rect 49374 233746 50048 233796
rect 47853 233744 50048 233746
rect 47853 233688 47858 233744
rect 47914 233736 50048 233744
rect 47914 233688 49434 233736
rect 47853 233686 49434 233688
rect 47853 233683 47919 233686
rect 48037 232794 48103 232797
rect 49374 232794 50048 232844
rect 48037 232792 50048 232794
rect 48037 232736 48042 232792
rect 48098 232784 50048 232792
rect 48098 232736 49434 232784
rect 48037 232734 49434 232736
rect 48037 232731 48103 232734
rect 237373 232522 237439 232525
rect 240182 232522 240242 233080
rect 237373 232520 240242 232522
rect 237373 232464 237378 232520
rect 237434 232464 240242 232520
rect 237373 232462 240242 232464
rect 237373 232459 237439 232462
rect 580073 232386 580139 232389
rect 583520 232386 584960 232476
rect 580073 232384 584960 232386
rect 580073 232328 580078 232384
rect 580134 232328 584960 232384
rect 580073 232326 584960 232328
rect 580073 232323 580139 232326
rect 238661 232114 238727 232117
rect 240182 232114 240242 232264
rect 583520 232236 584960 232326
rect 238661 232112 240242 232114
rect 238661 232056 238666 232112
rect 238722 232056 240242 232112
rect 238661 232054 240242 232056
rect 238661 232051 238727 232054
rect 47761 231026 47827 231029
rect 49374 231026 50048 231076
rect 47761 231024 50048 231026
rect 47761 230968 47766 231024
rect 47822 231016 50048 231024
rect 47822 230968 49434 231016
rect 47761 230966 49434 230968
rect 47761 230963 47827 230966
rect 237373 230210 237439 230213
rect 237373 230208 240242 230210
rect 237373 230152 237378 230208
rect 237434 230152 240242 230208
rect 237373 230150 240242 230152
rect 237373 230147 237439 230150
rect 47669 229938 47735 229941
rect 49374 229938 50048 229988
rect 47669 229936 50048 229938
rect 47669 229880 47674 229936
rect 47730 229928 50048 229936
rect 47730 229880 49434 229928
rect 47669 229878 49434 229880
rect 47669 229875 47735 229878
rect 240182 229600 240242 230150
rect 49509 228220 49575 228223
rect 49509 228218 50048 228220
rect 49509 228162 49514 228218
rect 49570 228162 50048 228218
rect 49509 228160 50048 228162
rect 237465 228170 237531 228173
rect 240182 228170 240242 228728
rect 237465 228168 240242 228170
rect 49509 228157 49575 228160
rect -960 227884 480 228124
rect 237465 228112 237470 228168
rect 237526 228112 240242 228168
rect 237465 228110 240242 228112
rect 237465 228107 237531 228110
rect 237373 227762 237439 227765
rect 240182 227762 240242 227776
rect 237373 227760 240242 227762
rect 237373 227704 237378 227760
rect 237434 227704 240242 227760
rect 237373 227702 240242 227704
rect 237373 227699 237439 227702
rect 238017 225858 238083 225861
rect 238017 225856 240242 225858
rect 238017 225800 238022 225856
rect 238078 225800 240242 225856
rect 238017 225798 240242 225800
rect 238017 225795 238083 225798
rect 240182 225248 240242 225798
rect 237373 223682 237439 223685
rect 240182 223682 240242 224240
rect 237373 223680 240242 223682
rect 237373 223624 237378 223680
rect 237434 223624 240242 223680
rect 237373 223622 240242 223624
rect 237373 223619 237439 223622
rect 237465 222866 237531 222869
rect 240182 222866 240242 223424
rect 237465 222864 240242 222866
rect 237465 222808 237470 222864
rect 237526 222808 240242 222864
rect 237465 222806 240242 222808
rect 237465 222803 237531 222806
rect 237373 222322 237439 222325
rect 240182 222322 240242 222608
rect 237373 222320 240242 222322
rect 237373 222264 237378 222320
rect 237434 222264 240242 222320
rect 237373 222262 240242 222264
rect 237373 222259 237439 222262
rect 237465 221642 237531 221645
rect 240182 221642 240242 221656
rect 237465 221640 240242 221642
rect 237465 221584 237470 221640
rect 237526 221584 240242 221640
rect 237465 221582 240242 221584
rect 237465 221579 237531 221582
rect 237373 221506 237439 221509
rect 237373 221504 240242 221506
rect 237373 221448 237378 221504
rect 237434 221448 240242 221504
rect 237373 221446 240242 221448
rect 237373 221443 237439 221446
rect 240182 220896 240242 221446
rect 237373 219602 237439 219605
rect 240182 219602 240242 219888
rect 237373 219600 240242 219602
rect 237373 219544 237378 219600
rect 237434 219544 240242 219600
rect 237373 219542 240242 219544
rect 237373 219539 237439 219542
rect 186588 219330 187250 219380
rect 189073 219330 189139 219333
rect 186588 219328 189139 219330
rect 186588 219320 189078 219328
rect 187190 219272 189078 219320
rect 189134 219272 189139 219328
rect 187190 219270 189139 219272
rect 189073 219267 189139 219270
rect 237465 218514 237531 218517
rect 240182 218514 240242 219072
rect 579797 219058 579863 219061
rect 583520 219058 584960 219148
rect 579797 219056 584960 219058
rect 579797 219000 579802 219056
rect 579858 219000 584960 219056
rect 579797 218998 584960 219000
rect 579797 218995 579863 218998
rect 583520 218908 584960 218998
rect 237465 218512 240242 218514
rect 237465 218456 237470 218512
rect 237526 218456 240242 218512
rect 237465 218454 240242 218456
rect 237465 218451 237531 218454
rect 237373 218106 237439 218109
rect 240182 218106 240242 218120
rect 237373 218104 240242 218106
rect 237373 218048 237378 218104
rect 237434 218048 240242 218104
rect 237373 218046 240242 218048
rect 237373 218043 237439 218046
rect 186588 217698 187250 217748
rect 189901 217698 189967 217701
rect 186588 217696 189967 217698
rect 186588 217688 189906 217696
rect 187190 217640 189906 217688
rect 189962 217640 189967 217696
rect 187190 217638 189967 217640
rect 189901 217635 189967 217638
rect 238518 216684 238524 216748
rect 238588 216746 238594 216748
rect 240182 216746 240242 217304
rect 238588 216686 240242 216746
rect 238588 216684 238594 216686
rect 237373 216474 237439 216477
rect 237373 216472 240242 216474
rect 237373 216416 237378 216472
rect 237434 216416 240242 216472
rect 237373 216414 240242 216416
rect 237373 216411 237439 216414
rect 240182 216408 240242 216414
rect 186588 216338 187250 216388
rect 189073 216338 189139 216341
rect 186588 216336 189139 216338
rect 186588 216328 189078 216336
rect 187190 216280 189078 216328
rect 189134 216280 189139 216336
rect 187190 216278 189139 216280
rect 189073 216275 189139 216278
rect 238017 215386 238083 215389
rect 240182 215386 240242 215536
rect 238017 215384 240242 215386
rect 238017 215328 238022 215384
rect 238078 215328 240242 215384
rect 238017 215326 240242 215328
rect 238017 215323 238083 215326
rect -960 214828 480 215068
rect 186588 214842 187250 214892
rect 190085 214842 190151 214845
rect 186588 214840 190151 214842
rect 186588 214832 190090 214840
rect 187190 214784 190090 214832
rect 190146 214784 190151 214840
rect 187190 214782 190151 214784
rect 190085 214779 190151 214782
rect 238293 214026 238359 214029
rect 240182 214026 240242 214584
rect 238293 214024 240242 214026
rect 238293 213968 238298 214024
rect 238354 213968 240242 214024
rect 238293 213966 240242 213968
rect 238293 213963 238359 213966
rect 186588 213618 187250 213668
rect 190269 213618 190335 213621
rect 186588 213616 190335 213618
rect 186588 213608 190274 213616
rect 187190 213560 190274 213608
rect 190330 213560 190335 213616
rect 187190 213558 190335 213560
rect 190269 213555 190335 213558
rect 237373 213482 237439 213485
rect 240182 213482 240242 213768
rect 237373 213480 240242 213482
rect 237373 213424 237378 213480
rect 237434 213424 240242 213480
rect 237373 213422 240242 213424
rect 237373 213419 237439 213422
rect 237465 212802 237531 212805
rect 240182 212802 240242 212952
rect 237465 212800 240242 212802
rect 237465 212744 237470 212800
rect 237526 212744 240242 212800
rect 237465 212742 240242 212744
rect 237465 212739 237531 212742
rect 237373 212394 237439 212397
rect 237373 212392 240242 212394
rect 237373 212336 237378 212392
rect 237434 212336 240242 212392
rect 237373 212334 240242 212336
rect 237373 212331 237439 212334
rect 240182 212056 240242 212334
rect 238477 211170 238543 211173
rect 240182 211170 240242 211184
rect 238477 211168 240242 211170
rect 238477 211112 238482 211168
rect 238538 211112 240242 211168
rect 238477 211110 240242 211112
rect 238477 211107 238543 211110
rect 49325 209946 49391 209949
rect 49742 209946 50048 209996
rect 49325 209944 50048 209946
rect 49325 209888 49330 209944
rect 49386 209936 50048 209944
rect 237465 209946 237531 209949
rect 240182 209946 240242 210232
rect 237465 209944 240242 209946
rect 49386 209888 49802 209936
rect 49325 209886 49802 209888
rect 237465 209888 237470 209944
rect 237526 209888 240242 209944
rect 237465 209886 240242 209888
rect 49325 209883 49391 209886
rect 237465 209883 237531 209886
rect 237373 209674 237439 209677
rect 237373 209672 240242 209674
rect 237373 209616 237378 209672
rect 237434 209616 240242 209672
rect 237373 209614 240242 209616
rect 237373 209611 237439 209614
rect 240182 209472 240242 209614
rect 237373 208450 237439 208453
rect 240182 208450 240242 208464
rect 237373 208448 240242 208450
rect 237373 208392 237378 208448
rect 237434 208392 240242 208448
rect 237373 208390 240242 208392
rect 237373 208387 237439 208390
rect 49601 208364 49667 208367
rect 49601 208362 50048 208364
rect 49601 208306 49606 208362
rect 49662 208306 50048 208362
rect 49601 208304 50048 208306
rect 237465 208314 237531 208317
rect 237465 208312 240242 208314
rect 49601 208301 49667 208304
rect 237465 208256 237470 208312
rect 237526 208256 240242 208312
rect 237465 208254 240242 208256
rect 237465 208251 237531 208254
rect 49417 208092 49483 208095
rect 49417 208090 50048 208092
rect 49417 208034 49422 208090
rect 49478 208034 50048 208090
rect 49417 208032 50048 208034
rect 49417 208029 49483 208032
rect 240182 207704 240242 208254
rect 237925 206138 237991 206141
rect 240182 206138 240242 206696
rect 237925 206136 240242 206138
rect 237925 206080 237930 206136
rect 237986 206080 240242 206136
rect 237925 206078 240242 206080
rect 237925 206075 237991 206078
rect 237465 205866 237531 205869
rect 240182 205866 240242 205880
rect 237465 205864 240242 205866
rect 237465 205808 237470 205864
rect 237526 205808 240242 205864
rect 237465 205806 240242 205808
rect 237465 205803 237531 205806
rect 187182 205668 187188 205732
rect 187252 205730 187258 205732
rect 187601 205730 187667 205733
rect 187252 205728 187667 205730
rect 187252 205672 187606 205728
rect 187662 205672 187667 205728
rect 187252 205670 187667 205672
rect 187252 205668 187258 205670
rect 187601 205667 187667 205670
rect 237373 205594 237439 205597
rect 237373 205592 240242 205594
rect 237373 205536 237378 205592
rect 237434 205536 240242 205592
rect 583520 205580 584960 205820
rect 237373 205534 240242 205536
rect 237373 205531 237439 205534
rect 240182 204984 240242 205534
rect 237373 203554 237439 203557
rect 240182 203554 240242 204112
rect 237373 203552 240242 203554
rect 237373 203496 237378 203552
rect 237434 203496 240242 203552
rect 237373 203494 240242 203496
rect 237373 203491 237439 203494
rect 237465 203010 237531 203013
rect 240182 203010 240242 203160
rect 237465 203008 240242 203010
rect 237465 202952 237470 203008
rect 237526 202952 240242 203008
rect 237465 202950 240242 202952
rect 237465 202947 237531 202950
rect 237373 202602 237439 202605
rect 237373 202600 240242 202602
rect 237373 202544 237378 202600
rect 237434 202544 240242 202600
rect 237373 202542 240242 202544
rect 237373 202539 237439 202542
rect 240182 202400 240242 202542
rect -960 201922 480 202012
rect 2773 201922 2839 201925
rect -960 201920 2839 201922
rect -960 201864 2778 201920
rect 2834 201864 2839 201920
rect -960 201862 2839 201864
rect -960 201772 480 201862
rect 2773 201859 2839 201862
rect 237373 201514 237439 201517
rect 240182 201514 240242 201528
rect 237373 201512 240242 201514
rect 237373 201456 237378 201512
rect 237434 201456 240242 201512
rect 237373 201454 240242 201456
rect 237373 201451 237439 201454
rect 237465 200154 237531 200157
rect 240182 200154 240242 200576
rect 237465 200152 240242 200154
rect 237465 200096 237470 200152
rect 237526 200096 240242 200152
rect 237465 200094 240242 200096
rect 237465 200091 237531 200094
rect 237373 200018 237439 200021
rect 237373 200016 240242 200018
rect 237373 199960 237378 200016
rect 237434 199960 240242 200016
rect 237373 199958 240242 199960
rect 237373 199955 237439 199958
rect 47945 199882 48011 199885
rect 238518 199882 238524 199884
rect 47945 199880 238524 199882
rect 47945 199824 47950 199880
rect 48006 199824 238524 199880
rect 47945 199822 238524 199824
rect 47945 199819 48011 199822
rect 238518 199820 238524 199822
rect 238588 199820 238594 199884
rect 240182 199816 240242 199958
rect 47853 199746 47919 199749
rect 234981 199746 235047 199749
rect 47853 199744 235047 199746
rect 47853 199688 47858 199744
rect 47914 199688 234986 199744
rect 235042 199688 235047 199744
rect 47853 199686 235047 199688
rect 47853 199683 47919 199686
rect 234981 199683 235047 199686
rect 48129 199610 48195 199613
rect 235165 199610 235231 199613
rect 48129 199608 235231 199610
rect 48129 199552 48134 199608
rect 48190 199552 235170 199608
rect 235226 199552 235231 199608
rect 48129 199550 235231 199552
rect 48129 199547 48195 199550
rect 235165 199547 235231 199550
rect 71865 199476 71931 199477
rect 77753 199476 77819 199477
rect 71814 199474 71820 199476
rect 71774 199414 71820 199474
rect 71884 199472 71931 199476
rect 77702 199474 77708 199476
rect 71926 199416 71931 199472
rect 71814 199412 71820 199414
rect 71884 199412 71931 199416
rect 77662 199414 77708 199474
rect 77772 199472 77819 199476
rect 77814 199416 77819 199472
rect 77702 199412 77708 199414
rect 77772 199412 77819 199416
rect 71865 199411 71931 199412
rect 77753 199411 77819 199412
rect 81341 199476 81407 199477
rect 82537 199476 82603 199477
rect 83457 199476 83523 199477
rect 86217 199476 86283 199477
rect 103697 199476 103763 199477
rect 150985 199476 151051 199477
rect 81341 199472 81388 199476
rect 81452 199474 81458 199476
rect 82486 199474 82492 199476
rect 81341 199416 81346 199472
rect 81341 199412 81388 199416
rect 81452 199414 81498 199474
rect 82446 199414 82492 199474
rect 82556 199472 82603 199476
rect 83406 199474 83412 199476
rect 82598 199416 82603 199472
rect 81452 199412 81458 199414
rect 82486 199412 82492 199414
rect 82556 199412 82603 199416
rect 83366 199414 83412 199474
rect 83476 199472 83523 199476
rect 86166 199474 86172 199476
rect 83518 199416 83523 199472
rect 83406 199412 83412 199414
rect 83476 199412 83523 199416
rect 86126 199414 86172 199474
rect 86236 199472 86283 199476
rect 103646 199474 103652 199476
rect 86278 199416 86283 199472
rect 86166 199412 86172 199414
rect 86236 199412 86283 199416
rect 103606 199414 103652 199474
rect 103716 199472 103763 199476
rect 150934 199474 150940 199476
rect 103758 199416 103763 199472
rect 103646 199412 103652 199414
rect 103716 199412 103763 199416
rect 150894 199414 150940 199474
rect 151004 199472 151051 199476
rect 151046 199416 151051 199472
rect 150934 199412 150940 199414
rect 151004 199412 151051 199416
rect 81341 199411 81407 199412
rect 82537 199411 82603 199412
rect 83457 199411 83523 199412
rect 86217 199411 86283 199412
rect 103697 199411 103763 199412
rect 150985 199411 151051 199412
rect 128353 199338 128419 199341
rect 237966 199338 237972 199340
rect 128353 199336 237972 199338
rect 128353 199280 128358 199336
rect 128414 199280 237972 199336
rect 128353 199278 237972 199280
rect 128353 199275 128419 199278
rect 237966 199276 237972 199278
rect 238036 199276 238042 199340
rect 47669 199066 47735 199069
rect 47669 199064 240242 199066
rect 47669 199008 47674 199064
rect 47730 199008 240242 199064
rect 47669 199006 240242 199008
rect 47669 199003 47735 199006
rect 103278 198868 103284 198932
rect 103348 198930 103354 198932
rect 186814 198930 186820 198932
rect 103348 198870 186820 198930
rect 103348 198868 103354 198870
rect 186814 198868 186820 198870
rect 186884 198868 186890 198932
rect 240182 198864 240242 199006
rect 70577 198660 70643 198661
rect 76649 198660 76715 198661
rect 78857 198660 78923 198661
rect 80145 198660 80211 198661
rect 84561 198660 84627 198661
rect 88241 198660 88307 198661
rect 88609 198660 88675 198661
rect 91185 198660 91251 198661
rect 93577 198660 93643 198661
rect 93945 198660 94011 198661
rect 95969 198660 96035 198661
rect 98361 198660 98427 198661
rect 99833 198660 99899 198661
rect 100937 198660 101003 198661
rect 102225 198660 102291 198661
rect 106089 198660 106155 198661
rect 107009 198660 107075 198661
rect 108481 198660 108547 198661
rect 113633 198660 113699 198661
rect 120993 198660 121059 198661
rect 123569 198660 123635 198661
rect 128537 198660 128603 198661
rect 130929 198660 130995 198661
rect 136081 198660 136147 198661
rect 70526 198658 70532 198660
rect 70486 198598 70532 198658
rect 70596 198656 70643 198660
rect 76598 198658 76604 198660
rect 70638 198600 70643 198656
rect 70526 198596 70532 198598
rect 70596 198596 70643 198600
rect 76558 198598 76604 198658
rect 76668 198656 76715 198660
rect 78806 198658 78812 198660
rect 76710 198600 76715 198656
rect 76598 198596 76604 198598
rect 76668 198596 76715 198600
rect 78766 198598 78812 198658
rect 78876 198656 78923 198660
rect 80094 198658 80100 198660
rect 78918 198600 78923 198656
rect 78806 198596 78812 198598
rect 78876 198596 78923 198600
rect 80054 198598 80100 198658
rect 80164 198656 80211 198660
rect 84510 198658 84516 198660
rect 80206 198600 80211 198656
rect 80094 198596 80100 198598
rect 80164 198596 80211 198600
rect 84470 198598 84516 198658
rect 84580 198656 84627 198660
rect 88190 198658 88196 198660
rect 84622 198600 84627 198656
rect 84510 198596 84516 198598
rect 84580 198596 84627 198600
rect 88150 198598 88196 198658
rect 88260 198656 88307 198660
rect 88558 198658 88564 198660
rect 88302 198600 88307 198656
rect 88190 198596 88196 198598
rect 88260 198596 88307 198600
rect 88518 198598 88564 198658
rect 88628 198656 88675 198660
rect 91134 198658 91140 198660
rect 88670 198600 88675 198656
rect 88558 198596 88564 198598
rect 88628 198596 88675 198600
rect 91094 198598 91140 198658
rect 91204 198656 91251 198660
rect 93526 198658 93532 198660
rect 91246 198600 91251 198656
rect 91134 198596 91140 198598
rect 91204 198596 91251 198600
rect 93486 198598 93532 198658
rect 93596 198656 93643 198660
rect 93894 198658 93900 198660
rect 93638 198600 93643 198656
rect 93526 198596 93532 198598
rect 93596 198596 93643 198600
rect 93854 198598 93900 198658
rect 93964 198656 94011 198660
rect 95918 198658 95924 198660
rect 94006 198600 94011 198656
rect 93894 198596 93900 198598
rect 93964 198596 94011 198600
rect 95878 198598 95924 198658
rect 95988 198656 96035 198660
rect 98310 198658 98316 198660
rect 96030 198600 96035 198656
rect 95918 198596 95924 198598
rect 95988 198596 96035 198600
rect 98270 198598 98316 198658
rect 98380 198656 98427 198660
rect 99782 198658 99788 198660
rect 98422 198600 98427 198656
rect 98310 198596 98316 198598
rect 98380 198596 98427 198600
rect 99742 198598 99788 198658
rect 99852 198656 99899 198660
rect 100886 198658 100892 198660
rect 99894 198600 99899 198656
rect 99782 198596 99788 198598
rect 99852 198596 99899 198600
rect 100846 198598 100892 198658
rect 100956 198656 101003 198660
rect 102174 198658 102180 198660
rect 100998 198600 101003 198656
rect 100886 198596 100892 198598
rect 100956 198596 101003 198600
rect 102134 198598 102180 198658
rect 102244 198656 102291 198660
rect 106038 198658 106044 198660
rect 102286 198600 102291 198656
rect 102174 198596 102180 198598
rect 102244 198596 102291 198600
rect 105998 198598 106044 198658
rect 106108 198656 106155 198660
rect 106958 198658 106964 198660
rect 106150 198600 106155 198656
rect 106038 198596 106044 198598
rect 106108 198596 106155 198600
rect 106918 198598 106964 198658
rect 107028 198656 107075 198660
rect 108430 198658 108436 198660
rect 107070 198600 107075 198656
rect 106958 198596 106964 198598
rect 107028 198596 107075 198600
rect 108390 198598 108436 198658
rect 108500 198656 108547 198660
rect 113582 198658 113588 198660
rect 108542 198600 108547 198656
rect 108430 198596 108436 198598
rect 108500 198596 108547 198600
rect 113542 198598 113588 198658
rect 113652 198656 113699 198660
rect 120942 198658 120948 198660
rect 113694 198600 113699 198656
rect 113582 198596 113588 198598
rect 113652 198596 113699 198600
rect 120902 198598 120948 198658
rect 121012 198656 121059 198660
rect 123518 198658 123524 198660
rect 121054 198600 121059 198656
rect 120942 198596 120948 198598
rect 121012 198596 121059 198600
rect 123478 198598 123524 198658
rect 123588 198656 123635 198660
rect 128486 198658 128492 198660
rect 123630 198600 123635 198656
rect 123518 198596 123524 198598
rect 123588 198596 123635 198600
rect 128446 198598 128492 198658
rect 128556 198656 128603 198660
rect 130878 198658 130884 198660
rect 128598 198600 128603 198656
rect 128486 198596 128492 198598
rect 128556 198596 128603 198600
rect 130838 198598 130884 198658
rect 130948 198656 130995 198660
rect 136030 198658 136036 198660
rect 130990 198600 130995 198656
rect 130878 198596 130884 198598
rect 130948 198596 130995 198600
rect 135990 198598 136036 198658
rect 136100 198656 136147 198660
rect 136142 198600 136147 198656
rect 136030 198596 136036 198598
rect 136100 198596 136147 198600
rect 138606 198596 138612 198660
rect 138676 198658 138682 198660
rect 138749 198658 138815 198661
rect 143441 198660 143507 198661
rect 146017 198660 146083 198661
rect 148593 198660 148659 198661
rect 153377 198660 153443 198661
rect 173433 198660 173499 198661
rect 143390 198658 143396 198660
rect 138676 198656 138815 198658
rect 138676 198600 138754 198656
rect 138810 198600 138815 198656
rect 138676 198598 138815 198600
rect 143350 198598 143396 198658
rect 143460 198656 143507 198660
rect 145966 198658 145972 198660
rect 143502 198600 143507 198656
rect 138676 198596 138682 198598
rect 70577 198595 70643 198596
rect 76649 198595 76715 198596
rect 78857 198595 78923 198596
rect 80145 198595 80211 198596
rect 84561 198595 84627 198596
rect 88241 198595 88307 198596
rect 88609 198595 88675 198596
rect 91185 198595 91251 198596
rect 93577 198595 93643 198596
rect 93945 198595 94011 198596
rect 95969 198595 96035 198596
rect 98361 198595 98427 198596
rect 99833 198595 99899 198596
rect 100937 198595 101003 198596
rect 102225 198595 102291 198596
rect 106089 198595 106155 198596
rect 107009 198595 107075 198596
rect 108481 198595 108547 198596
rect 113633 198595 113699 198596
rect 120993 198595 121059 198596
rect 123569 198595 123635 198596
rect 128537 198595 128603 198596
rect 130929 198595 130995 198596
rect 136081 198595 136147 198596
rect 138749 198595 138815 198598
rect 143390 198596 143396 198598
rect 143460 198596 143507 198600
rect 145926 198598 145972 198658
rect 146036 198656 146083 198660
rect 148542 198658 148548 198660
rect 146078 198600 146083 198656
rect 145966 198596 145972 198598
rect 146036 198596 146083 198600
rect 148502 198598 148548 198658
rect 148612 198656 148659 198660
rect 153326 198658 153332 198660
rect 148654 198600 148659 198656
rect 148542 198596 148548 198598
rect 148612 198596 148659 198600
rect 153286 198598 153332 198658
rect 153396 198656 153443 198660
rect 173382 198658 173388 198660
rect 153438 198600 153443 198656
rect 153326 198596 153332 198598
rect 153396 198596 153443 198600
rect 173342 198598 173388 198658
rect 173452 198656 173499 198660
rect 173494 198600 173499 198656
rect 173382 198596 173388 198598
rect 173452 198596 173499 198600
rect 143441 198595 143507 198596
rect 146017 198595 146083 198596
rect 148593 198595 148659 198596
rect 153377 198595 153443 198596
rect 173433 198595 173499 198596
rect 85849 198524 85915 198525
rect 85798 198522 85804 198524
rect 85758 198462 85804 198522
rect 85868 198520 85915 198524
rect 85910 198464 85915 198520
rect 85798 198460 85804 198462
rect 85868 198460 85915 198464
rect 87086 198460 87092 198524
rect 87156 198522 87162 198524
rect 87413 198522 87479 198525
rect 87156 198520 87479 198522
rect 87156 198464 87418 198520
rect 87474 198464 87479 198520
rect 87156 198462 87479 198464
rect 87156 198460 87162 198462
rect 85849 198459 85915 198460
rect 87413 198459 87479 198462
rect 90766 198460 90772 198524
rect 90836 198522 90842 198524
rect 90909 198522 90975 198525
rect 90836 198520 90975 198522
rect 90836 198464 90914 198520
rect 90970 198464 90975 198520
rect 90836 198462 90975 198464
rect 90836 198460 90842 198462
rect 90909 198459 90975 198462
rect 96470 198460 96476 198524
rect 96540 198522 96546 198524
rect 187141 198522 187207 198525
rect 96540 198520 187207 198522
rect 96540 198464 187146 198520
rect 187202 198464 187207 198520
rect 96540 198462 187207 198464
rect 96540 198460 96546 198462
rect 187141 198459 187207 198462
rect 89529 198388 89595 198389
rect 92841 198388 92907 198389
rect 89478 198386 89484 198388
rect 89438 198326 89484 198386
rect 89548 198384 89595 198388
rect 92790 198386 92796 198388
rect 89590 198328 89595 198384
rect 89478 198324 89484 198326
rect 89548 198324 89595 198328
rect 92750 198326 92796 198386
rect 92860 198384 92907 198388
rect 92902 198328 92907 198384
rect 92790 198324 92796 198326
rect 92860 198324 92907 198328
rect 95366 198324 95372 198388
rect 95436 198386 95442 198388
rect 187325 198386 187391 198389
rect 95436 198384 187391 198386
rect 95436 198328 187330 198384
rect 187386 198328 187391 198384
rect 95436 198326 187391 198328
rect 95436 198324 95442 198326
rect 89529 198323 89595 198324
rect 92841 198323 92907 198324
rect 187325 198323 187391 198326
rect 67214 198188 67220 198252
rect 67284 198250 67290 198252
rect 67541 198250 67607 198253
rect 67284 198248 67607 198250
rect 67284 198192 67546 198248
rect 67602 198192 67607 198248
rect 67284 198190 67607 198192
rect 67284 198188 67290 198190
rect 67541 198187 67607 198190
rect 74206 198188 74212 198252
rect 74276 198250 74282 198252
rect 74349 198250 74415 198253
rect 74276 198248 74415 198250
rect 74276 198192 74354 198248
rect 74410 198192 74415 198248
rect 74276 198190 74415 198192
rect 74276 198188 74282 198190
rect 74349 198187 74415 198190
rect 91870 198188 91876 198252
rect 91940 198250 91946 198252
rect 92289 198250 92355 198253
rect 91940 198248 92355 198250
rect 91940 198192 92294 198248
rect 92350 198192 92355 198248
rect 91940 198190 92355 198192
rect 91940 198188 91946 198190
rect 92289 198187 92355 198190
rect 101254 198188 101260 198252
rect 101324 198250 101330 198252
rect 186998 198250 187004 198252
rect 101324 198190 187004 198250
rect 101324 198188 101330 198190
rect 186998 198188 187004 198190
rect 187068 198188 187074 198252
rect 75494 198052 75500 198116
rect 75564 198114 75570 198116
rect 75729 198114 75795 198117
rect 75564 198112 75795 198114
rect 75564 198056 75734 198112
rect 75790 198056 75795 198112
rect 75564 198054 75795 198056
rect 75564 198052 75570 198054
rect 75729 198051 75795 198054
rect 104382 198052 104388 198116
rect 104452 198114 104458 198116
rect 187182 198114 187188 198116
rect 104452 198054 187188 198114
rect 104452 198052 104458 198054
rect 187182 198052 187188 198054
rect 187252 198052 187258 198116
rect 83590 197916 83596 197980
rect 83660 197978 83666 197980
rect 83733 197978 83799 197981
rect 105905 197980 105971 197981
rect 111057 197980 111123 197981
rect 105854 197978 105860 197980
rect 83660 197976 83799 197978
rect 83660 197920 83738 197976
rect 83794 197920 83799 197976
rect 83660 197918 83799 197920
rect 105814 197918 105860 197978
rect 105924 197976 105971 197980
rect 111006 197978 111012 197980
rect 105966 197920 105971 197976
rect 83660 197916 83666 197918
rect 83733 197915 83799 197918
rect 105854 197916 105860 197918
rect 105924 197916 105971 197920
rect 110966 197918 111012 197978
rect 111076 197976 111123 197980
rect 111118 197920 111123 197976
rect 111006 197916 111012 197918
rect 111076 197916 111123 197920
rect 140998 197916 141004 197980
rect 141068 197978 141074 197980
rect 188470 197978 188476 197980
rect 141068 197918 188476 197978
rect 141068 197916 141074 197918
rect 188470 197916 188476 197918
rect 188540 197916 188546 197980
rect 237373 197978 237439 197981
rect 240182 197978 240242 197992
rect 237373 197976 240242 197978
rect 237373 197920 237378 197976
rect 237434 197920 240242 197976
rect 237373 197918 240242 197920
rect 105905 197915 105971 197916
rect 111057 197915 111123 197916
rect 237373 197915 237439 197918
rect 115974 197780 115980 197844
rect 116044 197842 116050 197844
rect 116209 197842 116275 197845
rect 118417 197844 118483 197845
rect 155953 197844 156019 197845
rect 173249 197844 173315 197845
rect 118366 197842 118372 197844
rect 116044 197840 116275 197842
rect 116044 197784 116214 197840
rect 116270 197784 116275 197840
rect 116044 197782 116275 197784
rect 118326 197782 118372 197842
rect 118436 197840 118483 197844
rect 155902 197842 155908 197844
rect 118478 197784 118483 197840
rect 116044 197780 116050 197782
rect 116209 197779 116275 197782
rect 118366 197780 118372 197782
rect 118436 197780 118483 197784
rect 155862 197782 155908 197842
rect 155972 197840 156019 197844
rect 173198 197842 173204 197844
rect 156014 197784 156019 197840
rect 155902 197780 155908 197782
rect 155972 197780 156019 197784
rect 173158 197782 173204 197842
rect 173268 197840 173315 197844
rect 173310 197784 173315 197840
rect 173198 197780 173204 197782
rect 173268 197780 173315 197784
rect 118417 197779 118483 197780
rect 155953 197779 156019 197780
rect 173249 197779 173315 197780
rect 125910 197644 125916 197708
rect 125980 197706 125986 197708
rect 126145 197706 126211 197709
rect 133505 197708 133571 197709
rect 133454 197706 133460 197708
rect 125980 197704 126211 197706
rect 125980 197648 126150 197704
rect 126206 197648 126211 197704
rect 125980 197646 126211 197648
rect 133414 197646 133460 197706
rect 133524 197704 133571 197708
rect 133566 197648 133571 197704
rect 125980 197644 125986 197646
rect 126145 197643 126211 197646
rect 133454 197644 133460 197646
rect 133524 197644 133571 197648
rect 133505 197643 133571 197644
rect 98678 197508 98684 197572
rect 98748 197570 98754 197572
rect 238150 197570 238156 197572
rect 98748 197510 238156 197570
rect 98748 197508 98754 197510
rect 238150 197508 238156 197510
rect 238220 197508 238226 197572
rect 66161 197436 66227 197437
rect 66110 197434 66116 197436
rect 66070 197374 66116 197434
rect 66180 197432 66227 197436
rect 66222 197376 66227 197432
rect 66110 197372 66116 197374
rect 66180 197372 66227 197376
rect 68318 197372 68324 197436
rect 68388 197434 68394 197436
rect 68921 197434 68987 197437
rect 68388 197432 68987 197434
rect 68388 197376 68926 197432
rect 68982 197376 68987 197432
rect 68388 197374 68987 197376
rect 68388 197372 68394 197374
rect 66161 197371 66227 197372
rect 68921 197371 68987 197374
rect 69606 197372 69612 197436
rect 69676 197434 69682 197436
rect 69841 197434 69907 197437
rect 69676 197432 69907 197434
rect 69676 197376 69846 197432
rect 69902 197376 69907 197432
rect 69676 197374 69907 197376
rect 69676 197372 69682 197374
rect 69841 197371 69907 197374
rect 73102 197372 73108 197436
rect 73172 197434 73178 197436
rect 74441 197434 74507 197437
rect 73172 197432 74507 197434
rect 73172 197376 74446 197432
rect 74502 197376 74507 197432
rect 73172 197374 74507 197376
rect 73172 197372 73178 197374
rect 74441 197371 74507 197374
rect 78254 197372 78260 197436
rect 78324 197434 78330 197436
rect 78581 197434 78647 197437
rect 78324 197432 78647 197434
rect 78324 197376 78586 197432
rect 78642 197376 78647 197432
rect 78324 197374 78647 197376
rect 78324 197372 78330 197374
rect 78581 197371 78647 197374
rect 80830 197372 80836 197436
rect 80900 197434 80906 197436
rect 81065 197434 81131 197437
rect 80900 197432 81131 197434
rect 80900 197376 81070 197432
rect 81126 197376 81131 197432
rect 80900 197374 81131 197376
rect 80900 197372 80906 197374
rect 81065 197371 81131 197374
rect 97574 197372 97580 197436
rect 97644 197372 97650 197436
rect 97582 197298 97642 197372
rect 237373 197298 237439 197301
rect 97582 197238 235642 197298
rect 108062 197100 108068 197164
rect 108132 197162 108138 197164
rect 235441 197162 235507 197165
rect 108132 197160 235507 197162
rect 108132 197104 235446 197160
rect 235502 197104 235507 197160
rect 108132 197102 235507 197104
rect 235582 197162 235642 197238
rect 237373 197296 240242 197298
rect 237373 197240 237378 197296
rect 237434 197240 240242 197296
rect 237373 197238 240242 197240
rect 237373 197235 237439 197238
rect 238334 197162 238340 197164
rect 235582 197102 238340 197162
rect 108132 197100 108138 197102
rect 235441 197099 235507 197102
rect 238334 197100 238340 197102
rect 238404 197100 238410 197164
rect 240182 197096 240242 197238
rect 109166 196964 109172 197028
rect 109236 197026 109242 197028
rect 235574 197026 235580 197028
rect 109236 196966 235580 197026
rect 109236 196964 109242 196966
rect 235574 196964 235580 196966
rect 235644 196964 235650 197028
rect 138749 196890 138815 196893
rect 188654 196890 188660 196892
rect 138749 196888 188660 196890
rect 138749 196832 138754 196888
rect 138810 196832 188660 196888
rect 138749 196830 188660 196832
rect 138749 196827 138815 196830
rect 188654 196828 188660 196830
rect 188724 196828 188730 196892
rect 143441 196754 143507 196757
rect 188286 196754 188292 196756
rect 143441 196752 188292 196754
rect 143441 196696 143446 196752
rect 143502 196696 188292 196752
rect 143441 196694 188292 196696
rect 143441 196691 143507 196694
rect 188286 196692 188292 196694
rect 188356 196692 188362 196756
rect 237465 196074 237531 196077
rect 240182 196074 240242 196224
rect 237465 196072 240242 196074
rect 237465 196016 237470 196072
rect 237526 196016 240242 196072
rect 237465 196014 240242 196016
rect 237465 196011 237531 196014
rect 237373 195938 237439 195941
rect 237373 195936 240242 195938
rect 237373 195880 237378 195936
rect 237434 195880 240242 195936
rect 237373 195878 240242 195880
rect 237373 195875 237439 195878
rect 240182 195328 240242 195878
rect 237373 194442 237439 194445
rect 240182 194442 240242 194456
rect 237373 194440 240242 194442
rect 237373 194384 237378 194440
rect 237434 194384 240242 194440
rect 237373 194382 240242 194384
rect 237373 194379 237439 194382
rect 237465 194170 237531 194173
rect 237465 194168 240242 194170
rect 237465 194112 237470 194168
rect 237526 194112 240242 194168
rect 237465 194110 240242 194112
rect 237465 194107 237531 194110
rect 240182 193560 240242 194110
rect 237373 192946 237439 192949
rect 237373 192944 240242 192946
rect 237373 192888 237378 192944
rect 237434 192888 240242 192944
rect 237373 192886 240242 192888
rect 237373 192883 237439 192886
rect 240182 192744 240242 192886
rect 579981 192538 580047 192541
rect 583520 192538 584960 192628
rect 579981 192536 584960 192538
rect 579981 192480 579986 192536
rect 580042 192480 584960 192536
rect 579981 192478 584960 192480
rect 579981 192475 580047 192478
rect 583520 192388 584960 192478
rect 237465 191722 237531 191725
rect 240182 191722 240242 191736
rect 237465 191720 240242 191722
rect 237465 191664 237470 191720
rect 237526 191664 240242 191720
rect 237465 191662 240242 191664
rect 237465 191659 237531 191662
rect 237373 191586 237439 191589
rect 237373 191584 240242 191586
rect 237373 191528 237378 191584
rect 237434 191528 240242 191584
rect 237373 191526 240242 191528
rect 237373 191523 237439 191526
rect 240182 190976 240242 191526
rect 237373 190362 237439 190365
rect 237373 190360 240242 190362
rect 237373 190304 237378 190360
rect 237434 190304 240242 190360
rect 237373 190302 240242 190304
rect 237373 190299 237439 190302
rect 240182 190160 240242 190302
rect 237465 189818 237531 189821
rect 237465 189816 240242 189818
rect 237465 189760 237470 189816
rect 237526 189760 240242 189816
rect 237465 189758 240242 189760
rect 237465 189755 237531 189758
rect 240182 189208 240242 189758
rect 237373 189002 237439 189005
rect 237373 189000 240242 189002
rect -960 188866 480 188956
rect 237373 188944 237378 189000
rect 237434 188944 240242 189000
rect 237373 188942 240242 188944
rect 237373 188939 237439 188942
rect 3877 188866 3943 188869
rect -960 188864 3943 188866
rect -960 188808 3882 188864
rect 3938 188808 3943 188864
rect -960 188806 3943 188808
rect -960 188716 480 188806
rect 3877 188803 3943 188806
rect 240182 188392 240242 188942
rect 237373 187642 237439 187645
rect 237373 187640 240242 187642
rect 237373 187584 237378 187640
rect 237434 187584 240242 187640
rect 237373 187582 240242 187584
rect 237373 187579 237439 187582
rect 240182 187440 240242 187582
rect 235390 187172 235396 187236
rect 235460 187234 235466 187236
rect 235460 187174 240242 187234
rect 235460 187172 235466 187174
rect 240182 186624 240242 187174
rect 237373 186282 237439 186285
rect 237373 186280 240242 186282
rect 237373 186224 237378 186280
rect 237434 186224 240242 186280
rect 237373 186222 240242 186224
rect 237373 186219 237439 186222
rect 240182 185672 240242 186222
rect 237373 184922 237439 184925
rect 237373 184920 240242 184922
rect 237373 184864 237378 184920
rect 237434 184864 240242 184920
rect 237373 184862 240242 184864
rect 237373 184859 237439 184862
rect 240182 184856 240242 184862
rect 237465 184514 237531 184517
rect 237465 184512 240242 184514
rect 237465 184456 237470 184512
rect 237526 184456 240242 184512
rect 237465 184454 240242 184456
rect 237465 184451 237531 184454
rect 240182 183904 240242 184454
rect 237373 183290 237439 183293
rect 237373 183288 240242 183290
rect 237373 183232 237378 183288
rect 237434 183232 240242 183288
rect 237373 183230 240242 183232
rect 237373 183227 237439 183230
rect 240182 183088 240242 183230
rect 237373 182066 237439 182069
rect 240182 182066 240242 182080
rect 237373 182064 240242 182066
rect 237373 182008 237378 182064
rect 237434 182008 240242 182064
rect 237373 182006 240242 182008
rect 237373 182003 237439 182006
rect 490414 182004 490420 182068
rect 490484 182066 490490 182068
rect 491518 182066 491524 182068
rect 490484 182006 491524 182066
rect 490484 182004 490490 182006
rect 491518 182004 491524 182006
rect 491588 182004 491594 182068
rect 237465 181930 237531 181933
rect 237465 181928 240242 181930
rect 237465 181872 237470 181928
rect 237526 181872 240242 181928
rect 237465 181870 240242 181872
rect 237465 181867 237531 181870
rect 240182 181320 240242 181870
rect 237557 180706 237623 180709
rect 237557 180704 240242 180706
rect 237557 180648 237562 180704
rect 237618 180648 240242 180704
rect 237557 180646 240242 180648
rect 237557 180643 237623 180646
rect 240182 180472 240242 180646
rect 339033 179618 339099 179621
rect 580390 179618 580396 179620
rect 339033 179616 580396 179618
rect 339033 179560 339038 179616
rect 339094 179560 580396 179616
rect 339033 179558 580396 179560
rect 339033 179555 339099 179558
rect 580390 179556 580396 179558
rect 580460 179556 580466 179620
rect 7557 179482 7623 179485
rect 407665 179482 407731 179485
rect 7557 179480 407731 179482
rect 7557 179424 7562 179480
rect 7618 179424 407670 179480
rect 407726 179424 407731 179480
rect 7557 179422 407731 179424
rect 7557 179419 7623 179422
rect 407665 179419 407731 179422
rect 492673 179482 492739 179485
rect 494094 179482 494100 179484
rect 492673 179480 494100 179482
rect 492673 179424 492678 179480
rect 492734 179424 494100 179480
rect 492673 179422 494100 179424
rect 492673 179419 492739 179422
rect 494094 179420 494100 179422
rect 494164 179420 494170 179484
rect 235206 179284 235212 179348
rect 235276 179346 235282 179348
rect 466637 179346 466703 179349
rect 235276 179344 466703 179346
rect 235276 179288 466642 179344
rect 466698 179288 466703 179344
rect 235276 179286 466703 179288
rect 235276 179284 235282 179286
rect 466637 179283 466703 179286
rect 233969 179210 234035 179213
rect 425053 179210 425119 179213
rect 233969 179208 425119 179210
rect 233969 179152 233974 179208
rect 234030 179152 425058 179208
rect 425114 179152 425119 179208
rect 233969 179150 425119 179152
rect 233969 179147 234035 179150
rect 425053 179147 425119 179150
rect 580165 179210 580231 179213
rect 583520 179210 584960 179300
rect 580165 179208 584960 179210
rect 580165 179152 580170 179208
rect 580226 179152 584960 179208
rect 580165 179150 584960 179152
rect 580165 179147 580231 179150
rect 239254 179012 239260 179076
rect 239324 179074 239330 179076
rect 418153 179074 418219 179077
rect 239324 179072 418219 179074
rect 239324 179016 418158 179072
rect 418214 179016 418219 179072
rect 583520 179060 584960 179150
rect 239324 179014 418219 179016
rect 239324 179012 239330 179014
rect 418153 179011 418219 179014
rect 239489 178938 239555 178941
rect 411253 178938 411319 178941
rect 239489 178936 411319 178938
rect 239489 178880 239494 178936
rect 239550 178880 411258 178936
rect 411314 178880 411319 178936
rect 239489 178878 411319 178880
rect 239489 178875 239555 178878
rect 411253 178875 411319 178878
rect 485037 178938 485103 178941
rect 490414 178938 490420 178940
rect 485037 178936 490420 178938
rect 485037 178880 485042 178936
rect 485098 178880 490420 178936
rect 485037 178878 490420 178880
rect 485037 178875 485103 178878
rect 490414 178876 490420 178878
rect 490484 178876 490490 178940
rect 352833 178802 352899 178805
rect 491334 178802 491340 178804
rect 352833 178800 491340 178802
rect 352833 178744 352838 178800
rect 352894 178744 491340 178800
rect 352833 178742 491340 178744
rect 352833 178739 352899 178742
rect 491334 178740 491340 178742
rect 491404 178740 491410 178804
rect 370313 178666 370379 178669
rect 492806 178666 492812 178668
rect 370313 178664 492812 178666
rect 370313 178608 370318 178664
rect 370374 178608 492812 178664
rect 370313 178606 492812 178608
rect 370313 178603 370379 178606
rect 492806 178604 492812 178606
rect 492876 178604 492882 178668
rect 366541 177986 366607 177989
rect 379973 177986 380039 177989
rect 366541 177984 380039 177986
rect 366541 177928 366546 177984
rect 366602 177928 379978 177984
rect 380034 177928 380039 177984
rect 366541 177926 380039 177928
rect 366541 177923 366607 177926
rect 379973 177923 380039 177926
rect 356329 177850 356395 177853
rect 580206 177850 580212 177852
rect 356329 177848 580212 177850
rect 356329 177792 356334 177848
rect 356390 177792 580212 177848
rect 356329 177790 580212 177792
rect 356329 177787 356395 177790
rect 580206 177788 580212 177790
rect 580276 177788 580282 177852
rect 238753 177714 238819 177717
rect 435449 177714 435515 177717
rect 238753 177712 435515 177714
rect 238753 177656 238758 177712
rect 238814 177656 435454 177712
rect 435510 177656 435515 177712
rect 238753 177654 435515 177656
rect 238753 177651 238819 177654
rect 435449 177651 435515 177654
rect 237373 177578 237439 177581
rect 400765 177578 400831 177581
rect 237373 177576 400831 177578
rect 237373 177520 237378 177576
rect 237434 177520 400770 177576
rect 400826 177520 400831 177576
rect 237373 177518 400831 177520
rect 237373 177515 237439 177518
rect 400765 177515 400831 177518
rect 191189 177442 191255 177445
rect 442349 177442 442415 177445
rect 191189 177440 442415 177442
rect 191189 177384 191194 177440
rect 191250 177384 442354 177440
rect 442410 177384 442415 177440
rect 191189 177382 442415 177384
rect 191189 177379 191255 177382
rect 442349 177379 442415 177382
rect 332041 177306 332107 177309
rect 367001 177306 367067 177309
rect 332041 177304 367067 177306
rect 332041 177248 332046 177304
rect 332102 177248 367006 177304
rect 367062 177248 367067 177304
rect 332041 177246 367067 177248
rect 332041 177243 332107 177246
rect 367001 177243 367067 177246
rect -960 175796 480 176036
rect 583520 165732 584960 165972
rect -960 162740 480 162980
rect 580165 152690 580231 152693
rect 583520 152690 584960 152780
rect 580165 152688 584960 152690
rect 580165 152632 580170 152688
rect 580226 152632 584960 152688
rect 580165 152630 584960 152632
rect 580165 152627 580231 152630
rect 583520 152540 584960 152630
rect -960 149834 480 149924
rect 3417 149834 3483 149837
rect -960 149832 3483 149834
rect -960 149776 3422 149832
rect 3478 149776 3483 149832
rect -960 149774 3483 149776
rect -960 149684 480 149774
rect 3417 149771 3483 149774
rect 580165 139362 580231 139365
rect 583520 139362 584960 139452
rect 580165 139360 584960 139362
rect 580165 139304 580170 139360
rect 580226 139304 584960 139360
rect 580165 139302 584960 139304
rect 580165 139299 580231 139302
rect 583520 139212 584960 139302
rect -960 136778 480 136868
rect 3325 136778 3391 136781
rect -960 136776 3391 136778
rect -960 136720 3330 136776
rect 3386 136720 3391 136776
rect -960 136718 3391 136720
rect -960 136628 480 136718
rect 3325 136715 3391 136718
rect 583520 125884 584960 126124
rect -960 123572 480 123812
rect 579797 112842 579863 112845
rect 583520 112842 584960 112932
rect 579797 112840 584960 112842
rect 579797 112784 579802 112840
rect 579858 112784 584960 112840
rect 579797 112782 584960 112784
rect 579797 112779 579863 112782
rect 583520 112692 584960 112782
rect -960 110516 480 110756
rect 580165 99514 580231 99517
rect 583520 99514 584960 99604
rect 580165 99512 584960 99514
rect 580165 99456 580170 99512
rect 580226 99456 584960 99512
rect 580165 99454 584960 99456
rect 580165 99451 580231 99454
rect 583520 99364 584960 99454
rect -960 97460 480 97700
rect 583520 86036 584960 86276
rect -960 84690 480 84780
rect 3141 84690 3207 84693
rect -960 84688 3207 84690
rect -960 84632 3146 84688
rect 3202 84632 3207 84688
rect -960 84630 3207 84632
rect -960 84540 480 84630
rect 3141 84627 3207 84630
rect 580165 72994 580231 72997
rect 583520 72994 584960 73084
rect 580165 72992 584960 72994
rect 580165 72936 580170 72992
rect 580226 72936 584960 72992
rect 580165 72934 584960 72936
rect 580165 72931 580231 72934
rect 583520 72844 584960 72934
rect -960 71484 480 71724
rect 580165 59666 580231 59669
rect 583520 59666 584960 59756
rect 580165 59664 584960 59666
rect 580165 59608 580170 59664
rect 580226 59608 584960 59664
rect 580165 59606 584960 59608
rect 580165 59603 580231 59606
rect 583520 59516 584960 59606
rect -960 58428 480 58668
rect 583520 46188 584960 46428
rect -960 45522 480 45612
rect 3417 45522 3483 45525
rect -960 45520 3483 45522
rect -960 45464 3422 45520
rect 3478 45464 3483 45520
rect -960 45462 3483 45464
rect -960 45372 480 45462
rect 3417 45459 3483 45462
rect 580165 33146 580231 33149
rect 583520 33146 584960 33236
rect 580165 33144 584960 33146
rect 580165 33088 580170 33144
rect 580226 33088 584960 33144
rect 580165 33086 584960 33088
rect 580165 33083 580231 33086
rect 583520 32996 584960 33086
rect -960 32316 480 32556
rect 583520 19668 584960 19908
rect -960 19260 480 19500
rect 580165 6626 580231 6629
rect 583520 6626 584960 6716
rect 580165 6624 584960 6626
rect -960 6490 480 6580
rect 580165 6568 580170 6624
rect 580226 6568 584960 6624
rect 580165 6566 584960 6568
rect 580165 6563 580231 6566
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect 583520 6476 584960 6566
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
<< via3 >>
rect 491340 700436 491404 700500
rect 239260 700300 239324 700364
rect 492812 700300 492876 700364
rect 580212 697172 580276 697236
rect 580396 683844 580460 683908
rect 490420 498748 490484 498812
rect 494100 488548 494164 488612
rect 86172 466108 86236 466172
rect 237972 466108 238036 466172
rect 88564 465972 88628 466036
rect 93532 465836 93596 465900
rect 81020 465700 81084 465764
rect 78812 465564 78876 465628
rect 108436 465428 108500 465492
rect 238524 465428 238588 465492
rect 106228 465292 106292 465356
rect 238340 465292 238404 465356
rect 91140 465216 91204 465220
rect 91140 465160 91190 465216
rect 91190 465160 91204 465216
rect 91140 465156 91204 465160
rect 96108 465216 96172 465220
rect 96108 465160 96158 465216
rect 96158 465160 96172 465216
rect 96108 465156 96172 465160
rect 98500 465216 98564 465220
rect 98500 465160 98550 465216
rect 98550 465160 98564 465216
rect 98500 465156 98564 465160
rect 101260 465156 101324 465220
rect 103652 465216 103716 465220
rect 103652 465160 103702 465216
rect 103702 465160 103716 465216
rect 103652 465156 103716 465160
rect 111012 465216 111076 465220
rect 111012 465160 111062 465216
rect 111062 465160 111076 465216
rect 111012 465156 111076 465160
rect 113772 465216 113836 465220
rect 113772 465160 113822 465216
rect 113822 465160 113836 465216
rect 113772 465156 113836 465160
rect 116164 465216 116228 465220
rect 116164 465160 116214 465216
rect 116214 465160 116228 465216
rect 116164 465156 116228 465160
rect 118556 465216 118620 465220
rect 118556 465160 118606 465216
rect 118606 465160 118620 465216
rect 118556 465156 118620 465160
rect 128676 465216 128740 465220
rect 128676 465160 128726 465216
rect 128726 465160 128740 465216
rect 128676 465156 128740 465160
rect 136036 465216 136100 465220
rect 136036 465160 136086 465216
rect 136086 465160 136100 465216
rect 136036 465156 136100 465160
rect 141004 465216 141068 465220
rect 141004 465160 141054 465216
rect 141054 465160 141068 465216
rect 141004 465156 141068 465160
rect 143580 465216 143644 465220
rect 143580 465160 143630 465216
rect 143630 465160 143644 465216
rect 143580 465156 143644 465160
rect 153332 465216 153396 465220
rect 153332 465160 153382 465216
rect 153382 465160 153396 465216
rect 153332 465156 153396 465160
rect 156092 465216 156156 465220
rect 156092 465160 156142 465216
rect 156142 465160 156156 465216
rect 156092 465156 156156 465160
rect 168420 465216 168484 465220
rect 168420 465160 168470 465216
rect 168470 465160 168484 465216
rect 168420 465156 168484 465160
rect 169708 465216 169772 465220
rect 169708 465160 169758 465216
rect 169758 465160 169772 465216
rect 169708 465156 169772 465160
rect 180932 465156 180996 465220
rect 131068 463992 131132 463996
rect 131068 463936 131118 463992
rect 131118 463936 131132 463992
rect 131068 463932 131132 463936
rect 83462 463720 83526 463724
rect 83462 463664 83518 463720
rect 83518 463664 83526 463720
rect 83462 463660 83526 463664
rect 120998 463720 121062 463724
rect 120998 463664 121054 463720
rect 121054 463664 121062 463720
rect 120998 463660 121062 463664
rect 123582 463720 123646 463724
rect 123582 463664 123630 463720
rect 123630 463664 123646 463720
rect 123582 463660 123646 463664
rect 125894 463660 125958 463724
rect 133510 463720 133574 463724
rect 133510 463664 133566 463720
rect 133566 463664 133574 463720
rect 133510 463660 133574 463664
rect 138406 463660 138470 463724
rect 146022 463720 146086 463724
rect 146022 463664 146078 463720
rect 146078 463664 146086 463720
rect 146022 463660 146086 463664
rect 148470 463720 148534 463724
rect 148470 463664 148506 463720
rect 148506 463664 148534 463720
rect 148470 463660 148534 463664
rect 151054 463720 151118 463724
rect 151054 463664 151082 463720
rect 151082 463664 151118 463720
rect 151054 463660 151118 463664
rect 238156 461484 238220 461548
rect 490420 435916 490484 435980
rect 491524 435916 491588 435980
rect 123446 379672 123510 379676
rect 123446 379616 123482 379672
rect 123482 379616 123510 379672
rect 123446 379612 123510 379616
rect 130926 379672 130990 379676
rect 130926 379616 130934 379672
rect 130934 379616 130990 379672
rect 130926 379612 130990 379616
rect 133510 379672 133574 379676
rect 133510 379616 133566 379672
rect 133566 379616 133574 379672
rect 133510 379612 133574 379616
rect 145886 379672 145950 379676
rect 145886 379616 145930 379672
rect 145930 379616 145950 379672
rect 145886 379612 145950 379616
rect 148470 379672 148534 379676
rect 148470 379616 148506 379672
rect 148506 379616 148534 379672
rect 148470 379612 148534 379616
rect 155950 379672 156014 379676
rect 155950 379616 155958 379672
rect 155958 379616 156014 379672
rect 155950 379612 156014 379616
rect 93934 379536 93998 379540
rect 93934 379480 93950 379536
rect 93950 379480 93998 379536
rect 93934 379476 93998 379480
rect 96382 379536 96446 379540
rect 96382 379480 96434 379536
rect 96434 379480 96446 379536
rect 96382 379476 96446 379480
rect 97606 379536 97670 379540
rect 97606 379480 97630 379536
rect 97630 379480 97670 379536
rect 97606 379476 97670 379480
rect 98694 379536 98758 379540
rect 98694 379480 98734 379536
rect 98734 379480 98758 379536
rect 98694 379476 98758 379480
rect 102230 379536 102294 379540
rect 102230 379480 102286 379536
rect 102286 379480 102294 379536
rect 102230 379476 102294 379480
rect 125916 379536 125980 379540
rect 125916 379480 125966 379536
rect 125966 379480 125980 379536
rect 125916 379476 125980 379480
rect 128492 379536 128556 379540
rect 128492 379480 128542 379536
rect 128542 379480 128556 379536
rect 128492 379476 128556 379480
rect 108068 379340 108132 379404
rect 150940 379264 151004 379268
rect 150940 379208 150990 379264
rect 150990 379208 151004 379264
rect 150940 379204 151004 379208
rect 67220 378116 67284 378180
rect 74212 378116 74276 378180
rect 77708 378116 77772 378180
rect 81204 378116 81268 378180
rect 91876 378116 91940 378180
rect 95924 378116 95988 378180
rect 99788 378116 99852 378180
rect 103284 378116 103348 378180
rect 103652 378116 103716 378180
rect 113588 378116 113652 378180
rect 120948 378116 121012 378180
rect 153332 378116 153396 378180
rect 73108 378040 73172 378044
rect 73108 377984 73158 378040
rect 73158 377984 73172 378040
rect 73108 377980 73172 377984
rect 92796 378040 92860 378044
rect 92796 377984 92846 378040
rect 92846 377984 92860 378040
rect 92796 377980 92860 377984
rect 95188 377980 95252 378044
rect 101260 378040 101324 378044
rect 101260 377984 101310 378040
rect 101310 377984 101324 378040
rect 101260 377980 101324 377984
rect 105860 378040 105924 378044
rect 105860 377984 105910 378040
rect 105910 377984 105924 378040
rect 105860 377980 105924 377984
rect 106964 377980 107028 378044
rect 109172 377980 109236 378044
rect 136036 378040 136100 378044
rect 136036 377984 136086 378040
rect 136086 377984 136100 378040
rect 136036 377980 136100 377984
rect 138612 377980 138676 378044
rect 141004 377980 141068 378044
rect 143396 378040 143460 378044
rect 143396 377984 143446 378040
rect 143446 377984 143460 378040
rect 143396 377980 143460 377984
rect 104388 377904 104452 377908
rect 104388 377848 104438 377904
rect 104438 377848 104452 377904
rect 104388 377844 104452 377848
rect 66116 377088 66180 377092
rect 66116 377032 66166 377088
rect 66166 377032 66180 377088
rect 66116 377028 66180 377032
rect 68324 377028 68388 377092
rect 69612 377028 69676 377092
rect 70532 377028 70596 377092
rect 71820 377028 71884 377092
rect 75500 377028 75564 377092
rect 76604 377028 76668 377092
rect 78260 377088 78324 377092
rect 78260 377032 78310 377088
rect 78310 377032 78324 377088
rect 78260 377028 78324 377032
rect 78812 377028 78876 377092
rect 80100 377028 80164 377092
rect 82492 377028 82556 377092
rect 83596 377028 83660 377092
rect 84516 377028 84580 377092
rect 85988 377028 86052 377092
rect 88012 377028 88076 377092
rect 89484 377088 89548 377092
rect 89484 377032 89534 377088
rect 89534 377032 89548 377088
rect 89484 377028 89548 377032
rect 90772 377028 90836 377092
rect 91140 377028 91204 377092
rect 93532 377028 93596 377092
rect 98316 377028 98380 377092
rect 101076 377028 101140 377092
rect 106044 377028 106108 377092
rect 108436 377028 108500 377092
rect 111012 377028 111076 377092
rect 115980 377028 116044 377092
rect 118372 377028 118436 377092
rect 173388 377028 173452 377092
rect 80836 376892 80900 376956
rect 83412 376892 83476 376956
rect 85804 376892 85868 376956
rect 87092 376892 87156 376956
rect 88564 376892 88628 376956
rect 173204 376892 173268 376956
rect 238524 356628 238588 356692
rect 238340 351868 238404 351932
rect 235212 345068 235276 345132
rect 238156 329700 238220 329764
rect 237972 315964 238036 316028
rect 235580 290396 235644 290460
rect 136036 286180 136100 286244
rect 138428 286180 138492 286244
rect 143580 286180 143644 286244
rect 169708 286180 169772 286244
rect 78812 286044 78876 286108
rect 235396 286044 235460 286108
rect 106228 285968 106292 285972
rect 106228 285912 106242 285968
rect 106242 285912 106292 285968
rect 106228 285908 106292 285912
rect 108436 285908 108500 285972
rect 120764 285908 120828 285972
rect 187188 285908 187252 285972
rect 81020 285772 81084 285836
rect 83412 285636 83476 285700
rect 86172 285636 86236 285700
rect 88564 285636 88628 285700
rect 91140 285636 91204 285700
rect 93532 285636 93596 285700
rect 96292 285636 96356 285700
rect 103836 285636 103900 285700
rect 114324 285636 114388 285700
rect 118556 285696 118620 285700
rect 118556 285640 118606 285696
rect 118606 285640 118620 285696
rect 118556 285636 118620 285640
rect 123524 285636 123588 285700
rect 125916 285636 125980 285700
rect 133460 285636 133524 285700
rect 141004 285636 141068 285700
rect 151124 285636 151188 285700
rect 154068 285636 154132 285700
rect 156092 285636 156156 285700
rect 168420 285636 168484 285700
rect 128676 285152 128740 285156
rect 128676 285096 128726 285152
rect 128726 285096 128740 285152
rect 128676 285092 128740 285096
rect 131068 285152 131132 285156
rect 131068 285096 131118 285152
rect 131118 285096 131132 285152
rect 131068 285092 131132 285096
rect 111012 285016 111076 285020
rect 111012 284960 111062 285016
rect 111062 284960 111076 285016
rect 111012 284956 111076 284960
rect 116164 285016 116228 285020
rect 116164 284960 116214 285016
rect 116214 284960 116228 285016
rect 116164 284956 116228 284960
rect 98500 284880 98564 284884
rect 98500 284824 98550 284880
rect 98550 284824 98564 284880
rect 98500 284820 98564 284824
rect 148548 284880 148612 284884
rect 148548 284824 148598 284880
rect 148598 284824 148612 284880
rect 148548 284820 148612 284824
rect 101260 284744 101324 284748
rect 101260 284688 101310 284744
rect 101310 284688 101324 284744
rect 101260 284684 101324 284688
rect 145972 284744 146036 284748
rect 145972 284688 146022 284744
rect 146022 284688 146036 284744
rect 145972 284684 146036 284688
rect 180748 284064 180812 284068
rect 180748 284008 180762 284064
rect 180762 284008 180812 284064
rect 180748 284004 180812 284008
rect 188292 278972 188356 279036
rect 186820 277476 186884 277540
rect 188476 276116 188540 276180
rect 188660 273396 188724 273460
rect 187004 271900 187068 271964
rect 237972 269860 238036 269924
rect 238156 267276 238220 267340
rect 238340 264148 238404 264212
rect 187188 255308 187252 255372
rect 238524 216684 238588 216748
rect 187188 205668 187252 205732
rect 238524 199820 238588 199884
rect 71820 199472 71884 199476
rect 71820 199416 71870 199472
rect 71870 199416 71884 199472
rect 71820 199412 71884 199416
rect 77708 199472 77772 199476
rect 77708 199416 77758 199472
rect 77758 199416 77772 199472
rect 77708 199412 77772 199416
rect 81388 199472 81452 199476
rect 81388 199416 81402 199472
rect 81402 199416 81452 199472
rect 81388 199412 81452 199416
rect 82492 199472 82556 199476
rect 82492 199416 82542 199472
rect 82542 199416 82556 199472
rect 82492 199412 82556 199416
rect 83412 199472 83476 199476
rect 83412 199416 83462 199472
rect 83462 199416 83476 199472
rect 83412 199412 83476 199416
rect 86172 199472 86236 199476
rect 86172 199416 86222 199472
rect 86222 199416 86236 199472
rect 86172 199412 86236 199416
rect 103652 199472 103716 199476
rect 103652 199416 103702 199472
rect 103702 199416 103716 199472
rect 103652 199412 103716 199416
rect 150940 199472 151004 199476
rect 150940 199416 150990 199472
rect 150990 199416 151004 199472
rect 150940 199412 151004 199416
rect 237972 199276 238036 199340
rect 103284 198868 103348 198932
rect 186820 198868 186884 198932
rect 70532 198656 70596 198660
rect 70532 198600 70582 198656
rect 70582 198600 70596 198656
rect 70532 198596 70596 198600
rect 76604 198656 76668 198660
rect 76604 198600 76654 198656
rect 76654 198600 76668 198656
rect 76604 198596 76668 198600
rect 78812 198656 78876 198660
rect 78812 198600 78862 198656
rect 78862 198600 78876 198656
rect 78812 198596 78876 198600
rect 80100 198656 80164 198660
rect 80100 198600 80150 198656
rect 80150 198600 80164 198656
rect 80100 198596 80164 198600
rect 84516 198656 84580 198660
rect 84516 198600 84566 198656
rect 84566 198600 84580 198656
rect 84516 198596 84580 198600
rect 88196 198656 88260 198660
rect 88196 198600 88246 198656
rect 88246 198600 88260 198656
rect 88196 198596 88260 198600
rect 88564 198656 88628 198660
rect 88564 198600 88614 198656
rect 88614 198600 88628 198656
rect 88564 198596 88628 198600
rect 91140 198656 91204 198660
rect 91140 198600 91190 198656
rect 91190 198600 91204 198656
rect 91140 198596 91204 198600
rect 93532 198656 93596 198660
rect 93532 198600 93582 198656
rect 93582 198600 93596 198656
rect 93532 198596 93596 198600
rect 93900 198656 93964 198660
rect 93900 198600 93950 198656
rect 93950 198600 93964 198656
rect 93900 198596 93964 198600
rect 95924 198656 95988 198660
rect 95924 198600 95974 198656
rect 95974 198600 95988 198656
rect 95924 198596 95988 198600
rect 98316 198656 98380 198660
rect 98316 198600 98366 198656
rect 98366 198600 98380 198656
rect 98316 198596 98380 198600
rect 99788 198656 99852 198660
rect 99788 198600 99838 198656
rect 99838 198600 99852 198656
rect 99788 198596 99852 198600
rect 100892 198656 100956 198660
rect 100892 198600 100942 198656
rect 100942 198600 100956 198656
rect 100892 198596 100956 198600
rect 102180 198656 102244 198660
rect 102180 198600 102230 198656
rect 102230 198600 102244 198656
rect 102180 198596 102244 198600
rect 106044 198656 106108 198660
rect 106044 198600 106094 198656
rect 106094 198600 106108 198656
rect 106044 198596 106108 198600
rect 106964 198656 107028 198660
rect 106964 198600 107014 198656
rect 107014 198600 107028 198656
rect 106964 198596 107028 198600
rect 108436 198656 108500 198660
rect 108436 198600 108486 198656
rect 108486 198600 108500 198656
rect 108436 198596 108500 198600
rect 113588 198656 113652 198660
rect 113588 198600 113638 198656
rect 113638 198600 113652 198656
rect 113588 198596 113652 198600
rect 120948 198656 121012 198660
rect 120948 198600 120998 198656
rect 120998 198600 121012 198656
rect 120948 198596 121012 198600
rect 123524 198656 123588 198660
rect 123524 198600 123574 198656
rect 123574 198600 123588 198656
rect 123524 198596 123588 198600
rect 128492 198656 128556 198660
rect 128492 198600 128542 198656
rect 128542 198600 128556 198656
rect 128492 198596 128556 198600
rect 130884 198656 130948 198660
rect 130884 198600 130934 198656
rect 130934 198600 130948 198656
rect 130884 198596 130948 198600
rect 136036 198656 136100 198660
rect 136036 198600 136086 198656
rect 136086 198600 136100 198656
rect 136036 198596 136100 198600
rect 138612 198596 138676 198660
rect 143396 198656 143460 198660
rect 143396 198600 143446 198656
rect 143446 198600 143460 198656
rect 143396 198596 143460 198600
rect 145972 198656 146036 198660
rect 145972 198600 146022 198656
rect 146022 198600 146036 198656
rect 145972 198596 146036 198600
rect 148548 198656 148612 198660
rect 148548 198600 148598 198656
rect 148598 198600 148612 198656
rect 148548 198596 148612 198600
rect 153332 198656 153396 198660
rect 153332 198600 153382 198656
rect 153382 198600 153396 198656
rect 153332 198596 153396 198600
rect 173388 198656 173452 198660
rect 173388 198600 173438 198656
rect 173438 198600 173452 198656
rect 173388 198596 173452 198600
rect 85804 198520 85868 198524
rect 85804 198464 85854 198520
rect 85854 198464 85868 198520
rect 85804 198460 85868 198464
rect 87092 198460 87156 198524
rect 90772 198460 90836 198524
rect 96476 198460 96540 198524
rect 89484 198384 89548 198388
rect 89484 198328 89534 198384
rect 89534 198328 89548 198384
rect 89484 198324 89548 198328
rect 92796 198384 92860 198388
rect 92796 198328 92846 198384
rect 92846 198328 92860 198384
rect 92796 198324 92860 198328
rect 95372 198324 95436 198388
rect 67220 198188 67284 198252
rect 74212 198188 74276 198252
rect 91876 198188 91940 198252
rect 101260 198188 101324 198252
rect 187004 198188 187068 198252
rect 75500 198052 75564 198116
rect 104388 198052 104452 198116
rect 187188 198052 187252 198116
rect 83596 197916 83660 197980
rect 105860 197976 105924 197980
rect 105860 197920 105910 197976
rect 105910 197920 105924 197976
rect 105860 197916 105924 197920
rect 111012 197976 111076 197980
rect 111012 197920 111062 197976
rect 111062 197920 111076 197976
rect 111012 197916 111076 197920
rect 141004 197916 141068 197980
rect 188476 197916 188540 197980
rect 115980 197780 116044 197844
rect 118372 197840 118436 197844
rect 118372 197784 118422 197840
rect 118422 197784 118436 197840
rect 118372 197780 118436 197784
rect 155908 197840 155972 197844
rect 155908 197784 155958 197840
rect 155958 197784 155972 197840
rect 155908 197780 155972 197784
rect 173204 197840 173268 197844
rect 173204 197784 173254 197840
rect 173254 197784 173268 197840
rect 173204 197780 173268 197784
rect 125916 197644 125980 197708
rect 133460 197704 133524 197708
rect 133460 197648 133510 197704
rect 133510 197648 133524 197704
rect 133460 197644 133524 197648
rect 98684 197508 98748 197572
rect 238156 197508 238220 197572
rect 66116 197432 66180 197436
rect 66116 197376 66166 197432
rect 66166 197376 66180 197432
rect 66116 197372 66180 197376
rect 68324 197372 68388 197436
rect 69612 197372 69676 197436
rect 73108 197372 73172 197436
rect 78260 197372 78324 197436
rect 80836 197372 80900 197436
rect 97580 197372 97644 197436
rect 108068 197100 108132 197164
rect 238340 197100 238404 197164
rect 109172 196964 109236 197028
rect 235580 196964 235644 197028
rect 188660 196828 188724 196892
rect 188292 196692 188356 196756
rect 235396 187172 235460 187236
rect 490420 182004 490484 182068
rect 491524 182004 491588 182068
rect 580396 179556 580460 179620
rect 494100 179420 494164 179484
rect 235212 179284 235276 179348
rect 239260 179012 239324 179076
rect 490420 178876 490484 178940
rect 491340 178740 491404 178804
rect 492812 178604 492876 178668
rect 580212 177788 580276 177852
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 680614 -8106 711002
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 -8106 680614
rect -8726 680294 -8106 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 -8106 680294
rect -8726 644614 -8106 680058
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 -8106 644614
rect -8726 644294 -8106 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 -8106 644294
rect -8726 608614 -8106 644058
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 -8106 608614
rect -8726 608294 -8106 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 -8106 608294
rect -8726 572614 -8106 608058
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 -8106 572614
rect -8726 572294 -8106 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 -8106 572294
rect -8726 536614 -8106 572058
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 -8106 536614
rect -8726 536294 -8106 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 -8106 536294
rect -8726 500614 -8106 536058
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 -8106 500614
rect -8726 500294 -8106 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 -8106 500294
rect -8726 464614 -8106 500058
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 -8106 464614
rect -8726 464294 -8106 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 -8106 464294
rect -8726 428614 -8106 464058
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 -8106 428614
rect -8726 428294 -8106 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 -8106 428294
rect -8726 392614 -8106 428058
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 -8106 392614
rect -8726 392294 -8106 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 -8106 392294
rect -8726 356614 -8106 392058
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 -8106 356614
rect -8726 356294 -8106 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 -8106 356294
rect -8726 320614 -8106 356058
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 -8106 320614
rect -8726 320294 -8106 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 -8106 320294
rect -8726 284614 -8106 320058
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 -8106 284614
rect -8726 284294 -8106 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 -8106 284294
rect -8726 248614 -8106 284058
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 -8106 248614
rect -8726 248294 -8106 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 -8106 248294
rect -8726 212614 -8106 248058
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 -8106 212614
rect -8726 212294 -8106 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 -8106 212294
rect -8726 176614 -8106 212058
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 -8106 176614
rect -8726 176294 -8106 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 -8106 176294
rect -8726 140614 -8106 176058
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 -8106 140614
rect -8726 140294 -8106 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 -8106 140294
rect -8726 104614 -8106 140058
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 -8106 104614
rect -8726 104294 -8106 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 -8106 104294
rect -8726 68614 -8106 104058
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 -8106 68614
rect -8726 68294 -8106 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 -8106 68294
rect -8726 32614 -8106 68058
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 -8106 32614
rect -8726 32294 -8106 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 -8106 32294
rect -8726 -7066 -8106 32058
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 698614 -7146 710042
rect 12954 710598 13574 711590
rect 12954 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 13574 710598
rect 12954 710278 13574 710362
rect 12954 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 13574 710278
rect -7766 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 -7146 698614
rect -7766 698294 -7146 698378
rect -7766 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 -7146 698294
rect -7766 662614 -7146 698058
rect -7766 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 -7146 662614
rect -7766 662294 -7146 662378
rect -7766 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 -7146 662294
rect -7766 626614 -7146 662058
rect -7766 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 -7146 626614
rect -7766 626294 -7146 626378
rect -7766 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 -7146 626294
rect -7766 590614 -7146 626058
rect -7766 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 -7146 590614
rect -7766 590294 -7146 590378
rect -7766 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 -7146 590294
rect -7766 554614 -7146 590058
rect -7766 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 -7146 554614
rect -7766 554294 -7146 554378
rect -7766 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 -7146 554294
rect -7766 518614 -7146 554058
rect -7766 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 -7146 518614
rect -7766 518294 -7146 518378
rect -7766 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 -7146 518294
rect -7766 482614 -7146 518058
rect -7766 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 -7146 482614
rect -7766 482294 -7146 482378
rect -7766 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 -7146 482294
rect -7766 446614 -7146 482058
rect -7766 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 -7146 446614
rect -7766 446294 -7146 446378
rect -7766 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 -7146 446294
rect -7766 410614 -7146 446058
rect -7766 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 -7146 410614
rect -7766 410294 -7146 410378
rect -7766 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 -7146 410294
rect -7766 374614 -7146 410058
rect -7766 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 -7146 374614
rect -7766 374294 -7146 374378
rect -7766 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 -7146 374294
rect -7766 338614 -7146 374058
rect -7766 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 -7146 338614
rect -7766 338294 -7146 338378
rect -7766 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 -7146 338294
rect -7766 302614 -7146 338058
rect -7766 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 -7146 302614
rect -7766 302294 -7146 302378
rect -7766 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 -7146 302294
rect -7766 266614 -7146 302058
rect -7766 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 -7146 266614
rect -7766 266294 -7146 266378
rect -7766 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 -7146 266294
rect -7766 230614 -7146 266058
rect -7766 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 -7146 230614
rect -7766 230294 -7146 230378
rect -7766 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 -7146 230294
rect -7766 194614 -7146 230058
rect -7766 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 -7146 194614
rect -7766 194294 -7146 194378
rect -7766 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 -7146 194294
rect -7766 158614 -7146 194058
rect -7766 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 -7146 158614
rect -7766 158294 -7146 158378
rect -7766 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 -7146 158294
rect -7766 122614 -7146 158058
rect -7766 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 -7146 122614
rect -7766 122294 -7146 122378
rect -7766 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 -7146 122294
rect -7766 86614 -7146 122058
rect -7766 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 -7146 86614
rect -7766 86294 -7146 86378
rect -7766 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 -7146 86294
rect -7766 50614 -7146 86058
rect -7766 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 -7146 50614
rect -7766 50294 -7146 50378
rect -7766 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 -7146 50294
rect -7766 14614 -7146 50058
rect -7766 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 -7146 14614
rect -7766 14294 -7146 14378
rect -7766 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 -7146 14294
rect -7766 -6106 -7146 14058
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 676894 -6186 709082
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 -6186 676894
rect -6806 676574 -6186 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 -6186 676574
rect -6806 640894 -6186 676338
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 -6186 640894
rect -6806 640574 -6186 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 -6186 640574
rect -6806 604894 -6186 640338
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 -6186 604894
rect -6806 604574 -6186 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 -6186 604574
rect -6806 568894 -6186 604338
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 -6186 568894
rect -6806 568574 -6186 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 -6186 568574
rect -6806 532894 -6186 568338
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 -6186 532894
rect -6806 532574 -6186 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 -6186 532574
rect -6806 496894 -6186 532338
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 -6186 496894
rect -6806 496574 -6186 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 -6186 496574
rect -6806 460894 -6186 496338
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 -6186 460894
rect -6806 460574 -6186 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 -6186 460574
rect -6806 424894 -6186 460338
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 -6186 424894
rect -6806 424574 -6186 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 -6186 424574
rect -6806 388894 -6186 424338
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 -6186 388894
rect -6806 388574 -6186 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 -6186 388574
rect -6806 352894 -6186 388338
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 -6186 352894
rect -6806 352574 -6186 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 -6186 352574
rect -6806 316894 -6186 352338
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 -6186 316894
rect -6806 316574 -6186 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 -6186 316574
rect -6806 280894 -6186 316338
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 -6186 280894
rect -6806 280574 -6186 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 -6186 280574
rect -6806 244894 -6186 280338
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 -6186 244894
rect -6806 244574 -6186 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 -6186 244574
rect -6806 208894 -6186 244338
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 -6186 208894
rect -6806 208574 -6186 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 -6186 208574
rect -6806 172894 -6186 208338
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 -6186 172894
rect -6806 172574 -6186 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 -6186 172574
rect -6806 136894 -6186 172338
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 -6186 136894
rect -6806 136574 -6186 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 -6186 136574
rect -6806 100894 -6186 136338
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 -6186 100894
rect -6806 100574 -6186 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 -6186 100574
rect -6806 64894 -6186 100338
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 -6186 64894
rect -6806 64574 -6186 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 -6186 64574
rect -6806 28894 -6186 64338
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 -6186 28894
rect -6806 28574 -6186 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 -6186 28574
rect -6806 -5146 -6186 28338
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 694894 -5226 708122
rect 9234 708678 9854 709670
rect 9234 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 9854 708678
rect 9234 708358 9854 708442
rect 9234 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 9854 708358
rect -5846 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 -5226 694894
rect -5846 694574 -5226 694658
rect -5846 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 -5226 694574
rect -5846 658894 -5226 694338
rect -5846 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 -5226 658894
rect -5846 658574 -5226 658658
rect -5846 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 -5226 658574
rect -5846 622894 -5226 658338
rect -5846 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 -5226 622894
rect -5846 622574 -5226 622658
rect -5846 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 -5226 622574
rect -5846 586894 -5226 622338
rect -5846 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 -5226 586894
rect -5846 586574 -5226 586658
rect -5846 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 -5226 586574
rect -5846 550894 -5226 586338
rect -5846 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 -5226 550894
rect -5846 550574 -5226 550658
rect -5846 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 -5226 550574
rect -5846 514894 -5226 550338
rect -5846 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 -5226 514894
rect -5846 514574 -5226 514658
rect -5846 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 -5226 514574
rect -5846 478894 -5226 514338
rect -5846 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 -5226 478894
rect -5846 478574 -5226 478658
rect -5846 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 -5226 478574
rect -5846 442894 -5226 478338
rect -5846 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 -5226 442894
rect -5846 442574 -5226 442658
rect -5846 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 -5226 442574
rect -5846 406894 -5226 442338
rect -5846 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 -5226 406894
rect -5846 406574 -5226 406658
rect -5846 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 -5226 406574
rect -5846 370894 -5226 406338
rect -5846 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 -5226 370894
rect -5846 370574 -5226 370658
rect -5846 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 -5226 370574
rect -5846 334894 -5226 370338
rect -5846 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 -5226 334894
rect -5846 334574 -5226 334658
rect -5846 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 -5226 334574
rect -5846 298894 -5226 334338
rect -5846 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 -5226 298894
rect -5846 298574 -5226 298658
rect -5846 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 -5226 298574
rect -5846 262894 -5226 298338
rect -5846 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 -5226 262894
rect -5846 262574 -5226 262658
rect -5846 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 -5226 262574
rect -5846 226894 -5226 262338
rect -5846 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 -5226 226894
rect -5846 226574 -5226 226658
rect -5846 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 -5226 226574
rect -5846 190894 -5226 226338
rect -5846 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 -5226 190894
rect -5846 190574 -5226 190658
rect -5846 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 -5226 190574
rect -5846 154894 -5226 190338
rect -5846 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 -5226 154894
rect -5846 154574 -5226 154658
rect -5846 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 -5226 154574
rect -5846 118894 -5226 154338
rect -5846 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 -5226 118894
rect -5846 118574 -5226 118658
rect -5846 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 -5226 118574
rect -5846 82894 -5226 118338
rect -5846 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 -5226 82894
rect -5846 82574 -5226 82658
rect -5846 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 -5226 82574
rect -5846 46894 -5226 82338
rect -5846 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 -5226 46894
rect -5846 46574 -5226 46658
rect -5846 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 -5226 46574
rect -5846 10894 -5226 46338
rect -5846 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 -5226 10894
rect -5846 10574 -5226 10658
rect -5846 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 -5226 10574
rect -5846 -4186 -5226 10338
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 673174 -4266 707162
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 -4266 673174
rect -4886 672854 -4266 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 -4266 672854
rect -4886 637174 -4266 672618
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 -4266 637174
rect -4886 636854 -4266 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 -4266 636854
rect -4886 601174 -4266 636618
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 -4266 601174
rect -4886 600854 -4266 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 -4266 600854
rect -4886 565174 -4266 600618
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 -4266 565174
rect -4886 564854 -4266 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 -4266 564854
rect -4886 529174 -4266 564618
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 -4266 529174
rect -4886 528854 -4266 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 -4266 528854
rect -4886 493174 -4266 528618
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 -4266 493174
rect -4886 492854 -4266 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 -4266 492854
rect -4886 457174 -4266 492618
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 -4266 457174
rect -4886 456854 -4266 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 -4266 456854
rect -4886 421174 -4266 456618
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 -4266 421174
rect -4886 420854 -4266 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 -4266 420854
rect -4886 385174 -4266 420618
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 -4266 385174
rect -4886 384854 -4266 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 -4266 384854
rect -4886 349174 -4266 384618
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 -4266 349174
rect -4886 348854 -4266 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 -4266 348854
rect -4886 313174 -4266 348618
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 -4266 313174
rect -4886 312854 -4266 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 -4266 312854
rect -4886 277174 -4266 312618
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 -4266 277174
rect -4886 276854 -4266 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 -4266 276854
rect -4886 241174 -4266 276618
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 -4266 241174
rect -4886 240854 -4266 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 -4266 240854
rect -4886 205174 -4266 240618
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 -4266 205174
rect -4886 204854 -4266 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 -4266 204854
rect -4886 169174 -4266 204618
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 -4266 169174
rect -4886 168854 -4266 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 -4266 168854
rect -4886 133174 -4266 168618
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 -4266 133174
rect -4886 132854 -4266 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 -4266 132854
rect -4886 97174 -4266 132618
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 -4266 97174
rect -4886 96854 -4266 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 -4266 96854
rect -4886 61174 -4266 96618
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 -4266 61174
rect -4886 60854 -4266 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 -4266 60854
rect -4886 25174 -4266 60618
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 -4266 25174
rect -4886 24854 -4266 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 -4266 24854
rect -4886 -3226 -4266 24618
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 691174 -3306 706202
rect 5514 706758 6134 707750
rect 5514 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 6134 706758
rect 5514 706438 6134 706522
rect 5514 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 6134 706438
rect -3926 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 -3306 691174
rect -3926 690854 -3306 690938
rect -3926 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 -3306 690854
rect -3926 655174 -3306 690618
rect -3926 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 -3306 655174
rect -3926 654854 -3306 654938
rect -3926 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 -3306 654854
rect -3926 619174 -3306 654618
rect -3926 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 -3306 619174
rect -3926 618854 -3306 618938
rect -3926 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 -3306 618854
rect -3926 583174 -3306 618618
rect -3926 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 -3306 583174
rect -3926 582854 -3306 582938
rect -3926 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 -3306 582854
rect -3926 547174 -3306 582618
rect -3926 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 -3306 547174
rect -3926 546854 -3306 546938
rect -3926 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 -3306 546854
rect -3926 511174 -3306 546618
rect -3926 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 -3306 511174
rect -3926 510854 -3306 510938
rect -3926 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 -3306 510854
rect -3926 475174 -3306 510618
rect -3926 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 -3306 475174
rect -3926 474854 -3306 474938
rect -3926 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 -3306 474854
rect -3926 439174 -3306 474618
rect -3926 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 -3306 439174
rect -3926 438854 -3306 438938
rect -3926 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 -3306 438854
rect -3926 403174 -3306 438618
rect -3926 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 -3306 403174
rect -3926 402854 -3306 402938
rect -3926 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 -3306 402854
rect -3926 367174 -3306 402618
rect -3926 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 -3306 367174
rect -3926 366854 -3306 366938
rect -3926 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 -3306 366854
rect -3926 331174 -3306 366618
rect -3926 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 -3306 331174
rect -3926 330854 -3306 330938
rect -3926 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 -3306 330854
rect -3926 295174 -3306 330618
rect -3926 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 -3306 295174
rect -3926 294854 -3306 294938
rect -3926 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 -3306 294854
rect -3926 259174 -3306 294618
rect -3926 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 -3306 259174
rect -3926 258854 -3306 258938
rect -3926 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 -3306 258854
rect -3926 223174 -3306 258618
rect -3926 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 -3306 223174
rect -3926 222854 -3306 222938
rect -3926 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 -3306 222854
rect -3926 187174 -3306 222618
rect -3926 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 -3306 187174
rect -3926 186854 -3306 186938
rect -3926 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 -3306 186854
rect -3926 151174 -3306 186618
rect -3926 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 -3306 151174
rect -3926 150854 -3306 150938
rect -3926 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 -3306 150854
rect -3926 115174 -3306 150618
rect -3926 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 -3306 115174
rect -3926 114854 -3306 114938
rect -3926 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 -3306 114854
rect -3926 79174 -3306 114618
rect -3926 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 -3306 79174
rect -3926 78854 -3306 78938
rect -3926 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 -3306 78854
rect -3926 43174 -3306 78618
rect -3926 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 -3306 43174
rect -3926 42854 -3306 42938
rect -3926 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 -3306 42854
rect -3926 7174 -3306 42618
rect -3926 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 -3306 7174
rect -3926 6854 -3306 6938
rect -3926 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 -3306 6854
rect -3926 -2266 -3306 6618
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 669454 -2346 705242
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 -2346 669454
rect -2966 669134 -2346 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 -2346 669134
rect -2966 633454 -2346 668898
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 -2346 633454
rect -2966 633134 -2346 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 -2346 633134
rect -2966 597454 -2346 632898
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 -2346 597454
rect -2966 597134 -2346 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 -2346 597134
rect -2966 561454 -2346 596898
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 -2346 561454
rect -2966 561134 -2346 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 -2346 561134
rect -2966 525454 -2346 560898
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 -2346 525454
rect -2966 525134 -2346 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 -2346 525134
rect -2966 489454 -2346 524898
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 -2346 489454
rect -2966 489134 -2346 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 -2346 489134
rect -2966 453454 -2346 488898
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 -2346 453454
rect -2966 453134 -2346 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 -2346 453134
rect -2966 417454 -2346 452898
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 -2346 417454
rect -2966 417134 -2346 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 -2346 417134
rect -2966 381454 -2346 416898
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 -2346 381454
rect -2966 381134 -2346 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 -2346 381134
rect -2966 345454 -2346 380898
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 -2346 345454
rect -2966 345134 -2346 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 -2346 345134
rect -2966 309454 -2346 344898
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 -2346 309454
rect -2966 309134 -2346 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 -2346 309134
rect -2966 273454 -2346 308898
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 -2346 273454
rect -2966 273134 -2346 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 -2346 273134
rect -2966 237454 -2346 272898
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 -2346 237454
rect -2966 237134 -2346 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 -2346 237134
rect -2966 201454 -2346 236898
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 -2346 201454
rect -2966 201134 -2346 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 -2346 201134
rect -2966 165454 -2346 200898
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 -2346 165454
rect -2966 165134 -2346 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 -2346 165134
rect -2966 129454 -2346 164898
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 -2346 129454
rect -2966 129134 -2346 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 -2346 129134
rect -2966 93454 -2346 128898
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 -2346 93454
rect -2966 93134 -2346 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 -2346 93134
rect -2966 57454 -2346 92898
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 -2346 57454
rect -2966 57134 -2346 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 -2346 57134
rect -2966 21454 -2346 56898
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 -2346 21454
rect -2966 21134 -2346 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 -2346 21134
rect -2966 -1306 -2346 20898
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 705830
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 1794 -1894 2414 -902
rect 5514 691174 6134 706202
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect 5514 -2266 6134 6618
rect 5514 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 6134 -2266
rect 5514 -2586 6134 -2502
rect 5514 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 6134 -2586
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect 5514 -3814 6134 -2822
rect 9234 694894 9854 708122
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 658894 9854 694338
rect 9234 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 9854 658894
rect 9234 658574 9854 658658
rect 9234 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 9854 658574
rect 9234 622894 9854 658338
rect 9234 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 9854 622894
rect 9234 622574 9854 622658
rect 9234 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 9854 622574
rect 9234 586894 9854 622338
rect 9234 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 9854 586894
rect 9234 586574 9854 586658
rect 9234 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 9854 586574
rect 9234 550894 9854 586338
rect 9234 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 9854 550894
rect 9234 550574 9854 550658
rect 9234 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 9854 550574
rect 9234 514894 9854 550338
rect 9234 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 9854 514894
rect 9234 514574 9854 514658
rect 9234 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 9854 514574
rect 9234 478894 9854 514338
rect 9234 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 9854 478894
rect 9234 478574 9854 478658
rect 9234 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 9854 478574
rect 9234 442894 9854 478338
rect 9234 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 9854 442894
rect 9234 442574 9854 442658
rect 9234 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 9854 442574
rect 9234 406894 9854 442338
rect 9234 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 9854 406894
rect 9234 406574 9854 406658
rect 9234 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 9854 406574
rect 9234 370894 9854 406338
rect 9234 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 9854 370894
rect 9234 370574 9854 370658
rect 9234 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 9854 370574
rect 9234 334894 9854 370338
rect 9234 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 9854 334894
rect 9234 334574 9854 334658
rect 9234 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 9854 334574
rect 9234 298894 9854 334338
rect 9234 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 9854 298894
rect 9234 298574 9854 298658
rect 9234 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 9854 298574
rect 9234 262894 9854 298338
rect 9234 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 9854 262894
rect 9234 262574 9854 262658
rect 9234 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 9854 262574
rect 9234 226894 9854 262338
rect 9234 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 9854 226894
rect 9234 226574 9854 226658
rect 9234 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 9854 226574
rect 9234 190894 9854 226338
rect 9234 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 9854 190894
rect 9234 190574 9854 190658
rect 9234 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 9854 190574
rect 9234 154894 9854 190338
rect 9234 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 9854 154894
rect 9234 154574 9854 154658
rect 9234 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 9854 154574
rect 9234 118894 9854 154338
rect 9234 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 9854 118894
rect 9234 118574 9854 118658
rect 9234 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 9854 118574
rect 9234 82894 9854 118338
rect 9234 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 9854 82894
rect 9234 82574 9854 82658
rect 9234 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 9854 82574
rect 9234 46894 9854 82338
rect 9234 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 9854 46894
rect 9234 46574 9854 46658
rect 9234 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 9854 46574
rect 9234 10894 9854 46338
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect 9234 -4186 9854 10338
rect 9234 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 9854 -4186
rect 9234 -4506 9854 -4422
rect 9234 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 9854 -4506
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect 9234 -5734 9854 -4742
rect 12954 698614 13574 710042
rect 30954 711558 31574 711590
rect 30954 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 31574 711558
rect 30954 711238 31574 711322
rect 30954 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 31574 711238
rect 27234 709638 27854 709670
rect 27234 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 27854 709638
rect 27234 709318 27854 709402
rect 27234 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 27854 709318
rect 23514 707718 24134 707750
rect 23514 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 24134 707718
rect 23514 707398 24134 707482
rect 23514 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 24134 707398
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 662614 13574 698058
rect 12954 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 13574 662614
rect 12954 662294 13574 662378
rect 12954 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 13574 662294
rect 12954 626614 13574 662058
rect 12954 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 13574 626614
rect 12954 626294 13574 626378
rect 12954 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 13574 626294
rect 12954 590614 13574 626058
rect 12954 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 13574 590614
rect 12954 590294 13574 590378
rect 12954 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 13574 590294
rect 12954 554614 13574 590058
rect 12954 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 13574 554614
rect 12954 554294 13574 554378
rect 12954 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 13574 554294
rect 12954 518614 13574 554058
rect 12954 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 13574 518614
rect 12954 518294 13574 518378
rect 12954 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 13574 518294
rect 12954 482614 13574 518058
rect 12954 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 13574 482614
rect 12954 482294 13574 482378
rect 12954 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 13574 482294
rect 12954 446614 13574 482058
rect 12954 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 13574 446614
rect 12954 446294 13574 446378
rect 12954 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 13574 446294
rect 12954 410614 13574 446058
rect 12954 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 13574 410614
rect 12954 410294 13574 410378
rect 12954 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 13574 410294
rect 12954 374614 13574 410058
rect 12954 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 13574 374614
rect 12954 374294 13574 374378
rect 12954 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 13574 374294
rect 12954 338614 13574 374058
rect 12954 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 13574 338614
rect 12954 338294 13574 338378
rect 12954 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 13574 338294
rect 12954 302614 13574 338058
rect 12954 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 13574 302614
rect 12954 302294 13574 302378
rect 12954 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 13574 302294
rect 12954 266614 13574 302058
rect 12954 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 13574 266614
rect 12954 266294 13574 266378
rect 12954 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 13574 266294
rect 12954 230614 13574 266058
rect 12954 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 13574 230614
rect 12954 230294 13574 230378
rect 12954 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 13574 230294
rect 12954 194614 13574 230058
rect 12954 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 13574 194614
rect 12954 194294 13574 194378
rect 12954 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 13574 194294
rect 12954 158614 13574 194058
rect 12954 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 13574 158614
rect 12954 158294 13574 158378
rect 12954 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 13574 158294
rect 12954 122614 13574 158058
rect 12954 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 13574 122614
rect 12954 122294 13574 122378
rect 12954 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 13574 122294
rect 12954 86614 13574 122058
rect 12954 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 13574 86614
rect 12954 86294 13574 86378
rect 12954 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 13574 86294
rect 12954 50614 13574 86058
rect 12954 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 13574 50614
rect 12954 50294 13574 50378
rect 12954 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 13574 50294
rect 12954 14614 13574 50058
rect 12954 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 13574 14614
rect 12954 14294 13574 14378
rect 12954 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 13574 14294
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect 12954 -6106 13574 14058
rect 19794 705798 20414 705830
rect 19794 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 20414 705798
rect 19794 705478 20414 705562
rect 19794 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 20414 705478
rect 19794 669454 20414 705242
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -1306 20414 20898
rect 19794 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 20414 -1306
rect 19794 -1626 20414 -1542
rect 19794 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 20414 -1626
rect 19794 -1894 20414 -1862
rect 23514 673174 24134 707162
rect 23514 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 24134 673174
rect 23514 672854 24134 672938
rect 23514 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 24134 672854
rect 23514 637174 24134 672618
rect 23514 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 24134 637174
rect 23514 636854 24134 636938
rect 23514 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 24134 636854
rect 23514 601174 24134 636618
rect 23514 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 24134 601174
rect 23514 600854 24134 600938
rect 23514 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 24134 600854
rect 23514 565174 24134 600618
rect 23514 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 24134 565174
rect 23514 564854 24134 564938
rect 23514 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 24134 564854
rect 23514 529174 24134 564618
rect 23514 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 24134 529174
rect 23514 528854 24134 528938
rect 23514 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 24134 528854
rect 23514 493174 24134 528618
rect 23514 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 24134 493174
rect 23514 492854 24134 492938
rect 23514 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 24134 492854
rect 23514 457174 24134 492618
rect 23514 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 24134 457174
rect 23514 456854 24134 456938
rect 23514 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 24134 456854
rect 23514 421174 24134 456618
rect 23514 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 24134 421174
rect 23514 420854 24134 420938
rect 23514 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 24134 420854
rect 23514 385174 24134 420618
rect 23514 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 24134 385174
rect 23514 384854 24134 384938
rect 23514 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 24134 384854
rect 23514 349174 24134 384618
rect 23514 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 24134 349174
rect 23514 348854 24134 348938
rect 23514 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 24134 348854
rect 23514 313174 24134 348618
rect 23514 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 24134 313174
rect 23514 312854 24134 312938
rect 23514 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 24134 312854
rect 23514 277174 24134 312618
rect 23514 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 24134 277174
rect 23514 276854 24134 276938
rect 23514 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 24134 276854
rect 23514 241174 24134 276618
rect 23514 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 24134 241174
rect 23514 240854 24134 240938
rect 23514 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 24134 240854
rect 23514 205174 24134 240618
rect 23514 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 24134 205174
rect 23514 204854 24134 204938
rect 23514 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 24134 204854
rect 23514 169174 24134 204618
rect 23514 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 24134 169174
rect 23514 168854 24134 168938
rect 23514 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 24134 168854
rect 23514 133174 24134 168618
rect 23514 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 24134 133174
rect 23514 132854 24134 132938
rect 23514 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 24134 132854
rect 23514 97174 24134 132618
rect 23514 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 24134 97174
rect 23514 96854 24134 96938
rect 23514 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 24134 96854
rect 23514 61174 24134 96618
rect 23514 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 24134 61174
rect 23514 60854 24134 60938
rect 23514 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 24134 60854
rect 23514 25174 24134 60618
rect 23514 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 24134 25174
rect 23514 24854 24134 24938
rect 23514 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 24134 24854
rect 23514 -3226 24134 24618
rect 23514 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 24134 -3226
rect 23514 -3546 24134 -3462
rect 23514 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 24134 -3546
rect 23514 -3814 24134 -3782
rect 27234 676894 27854 709082
rect 27234 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 27854 676894
rect 27234 676574 27854 676658
rect 27234 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 27854 676574
rect 27234 640894 27854 676338
rect 27234 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 27854 640894
rect 27234 640574 27854 640658
rect 27234 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 27854 640574
rect 27234 604894 27854 640338
rect 27234 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 27854 604894
rect 27234 604574 27854 604658
rect 27234 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 27854 604574
rect 27234 568894 27854 604338
rect 27234 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 27854 568894
rect 27234 568574 27854 568658
rect 27234 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 27854 568574
rect 27234 532894 27854 568338
rect 27234 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 27854 532894
rect 27234 532574 27854 532658
rect 27234 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 27854 532574
rect 27234 496894 27854 532338
rect 27234 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 27854 496894
rect 27234 496574 27854 496658
rect 27234 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 27854 496574
rect 27234 460894 27854 496338
rect 27234 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 27854 460894
rect 27234 460574 27854 460658
rect 27234 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 27854 460574
rect 27234 424894 27854 460338
rect 27234 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 27854 424894
rect 27234 424574 27854 424658
rect 27234 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 27854 424574
rect 27234 388894 27854 424338
rect 27234 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 27854 388894
rect 27234 388574 27854 388658
rect 27234 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 27854 388574
rect 27234 352894 27854 388338
rect 27234 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 27854 352894
rect 27234 352574 27854 352658
rect 27234 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 27854 352574
rect 27234 316894 27854 352338
rect 27234 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 27854 316894
rect 27234 316574 27854 316658
rect 27234 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 27854 316574
rect 27234 280894 27854 316338
rect 27234 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 27854 280894
rect 27234 280574 27854 280658
rect 27234 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 27854 280574
rect 27234 244894 27854 280338
rect 27234 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 27854 244894
rect 27234 244574 27854 244658
rect 27234 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 27854 244574
rect 27234 208894 27854 244338
rect 27234 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 27854 208894
rect 27234 208574 27854 208658
rect 27234 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 27854 208574
rect 27234 172894 27854 208338
rect 27234 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 27854 172894
rect 27234 172574 27854 172658
rect 27234 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 27854 172574
rect 27234 136894 27854 172338
rect 27234 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 27854 136894
rect 27234 136574 27854 136658
rect 27234 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 27854 136574
rect 27234 100894 27854 136338
rect 27234 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 27854 100894
rect 27234 100574 27854 100658
rect 27234 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 27854 100574
rect 27234 64894 27854 100338
rect 27234 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 27854 64894
rect 27234 64574 27854 64658
rect 27234 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 27854 64574
rect 27234 28894 27854 64338
rect 27234 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 27854 28894
rect 27234 28574 27854 28658
rect 27234 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 27854 28574
rect 27234 -5146 27854 28338
rect 27234 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 27854 -5146
rect 27234 -5466 27854 -5382
rect 27234 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 27854 -5466
rect 27234 -5734 27854 -5702
rect 30954 680614 31574 711002
rect 48954 710598 49574 711590
rect 48954 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 49574 710598
rect 48954 710278 49574 710362
rect 48954 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 49574 710278
rect 45234 708678 45854 709670
rect 45234 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 45854 708678
rect 45234 708358 45854 708442
rect 45234 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 45854 708358
rect 41514 706758 42134 707750
rect 41514 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 42134 706758
rect 41514 706438 42134 706522
rect 41514 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 42134 706438
rect 30954 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 31574 680614
rect 30954 680294 31574 680378
rect 30954 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 31574 680294
rect 30954 644614 31574 680058
rect 30954 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 31574 644614
rect 30954 644294 31574 644378
rect 30954 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 31574 644294
rect 30954 608614 31574 644058
rect 30954 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 31574 608614
rect 30954 608294 31574 608378
rect 30954 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 31574 608294
rect 30954 572614 31574 608058
rect 30954 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 31574 572614
rect 30954 572294 31574 572378
rect 30954 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 31574 572294
rect 30954 536614 31574 572058
rect 30954 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 31574 536614
rect 30954 536294 31574 536378
rect 30954 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 31574 536294
rect 30954 500614 31574 536058
rect 30954 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 31574 500614
rect 30954 500294 31574 500378
rect 30954 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 31574 500294
rect 30954 464614 31574 500058
rect 30954 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 31574 464614
rect 30954 464294 31574 464378
rect 30954 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 31574 464294
rect 30954 428614 31574 464058
rect 30954 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 31574 428614
rect 30954 428294 31574 428378
rect 30954 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 31574 428294
rect 30954 392614 31574 428058
rect 30954 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 31574 392614
rect 30954 392294 31574 392378
rect 30954 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 31574 392294
rect 30954 356614 31574 392058
rect 30954 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 31574 356614
rect 30954 356294 31574 356378
rect 30954 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 31574 356294
rect 30954 320614 31574 356058
rect 30954 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 31574 320614
rect 30954 320294 31574 320378
rect 30954 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 31574 320294
rect 30954 284614 31574 320058
rect 30954 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 31574 284614
rect 30954 284294 31574 284378
rect 30954 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 31574 284294
rect 30954 248614 31574 284058
rect 30954 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 31574 248614
rect 30954 248294 31574 248378
rect 30954 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 31574 248294
rect 30954 212614 31574 248058
rect 30954 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 31574 212614
rect 30954 212294 31574 212378
rect 30954 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 31574 212294
rect 30954 176614 31574 212058
rect 30954 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 31574 176614
rect 30954 176294 31574 176378
rect 30954 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 31574 176294
rect 30954 140614 31574 176058
rect 30954 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 31574 140614
rect 30954 140294 31574 140378
rect 30954 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 31574 140294
rect 30954 104614 31574 140058
rect 30954 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 31574 104614
rect 30954 104294 31574 104378
rect 30954 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 31574 104294
rect 30954 68614 31574 104058
rect 30954 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 31574 68614
rect 30954 68294 31574 68378
rect 30954 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 31574 68294
rect 30954 32614 31574 68058
rect 30954 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 31574 32614
rect 30954 32294 31574 32378
rect 30954 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 31574 32294
rect 12954 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 13574 -6106
rect 12954 -6426 13574 -6342
rect 12954 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 13574 -6426
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 12954 -7654 13574 -6662
rect 30954 -7066 31574 32058
rect 37794 704838 38414 705830
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -1894 38414 -902
rect 41514 691174 42134 706202
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 41514 655174 42134 690618
rect 41514 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 42134 655174
rect 41514 654854 42134 654938
rect 41514 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 42134 654854
rect 41514 619174 42134 654618
rect 41514 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 42134 619174
rect 41514 618854 42134 618938
rect 41514 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 42134 618854
rect 41514 583174 42134 618618
rect 41514 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 42134 583174
rect 41514 582854 42134 582938
rect 41514 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 42134 582854
rect 41514 547174 42134 582618
rect 41514 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 42134 547174
rect 41514 546854 42134 546938
rect 41514 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 42134 546854
rect 41514 511174 42134 546618
rect 41514 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 42134 511174
rect 41514 510854 42134 510938
rect 41514 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 42134 510854
rect 41514 475174 42134 510618
rect 41514 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 42134 475174
rect 41514 474854 42134 474938
rect 41514 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 42134 474854
rect 41514 439174 42134 474618
rect 41514 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 42134 439174
rect 41514 438854 42134 438938
rect 41514 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 42134 438854
rect 41514 403174 42134 438618
rect 41514 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 42134 403174
rect 41514 402854 42134 402938
rect 41514 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 42134 402854
rect 41514 367174 42134 402618
rect 41514 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 42134 367174
rect 41514 366854 42134 366938
rect 41514 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 42134 366854
rect 41514 331174 42134 366618
rect 41514 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 42134 331174
rect 41514 330854 42134 330938
rect 41514 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 42134 330854
rect 41514 295174 42134 330618
rect 41514 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 42134 295174
rect 41514 294854 42134 294938
rect 41514 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 42134 294854
rect 41514 259174 42134 294618
rect 41514 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 42134 259174
rect 41514 258854 42134 258938
rect 41514 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 42134 258854
rect 41514 223174 42134 258618
rect 41514 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 42134 223174
rect 41514 222854 42134 222938
rect 41514 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 42134 222854
rect 41514 187174 42134 222618
rect 41514 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 42134 187174
rect 41514 186854 42134 186938
rect 41514 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 42134 186854
rect 41514 151174 42134 186618
rect 41514 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 42134 151174
rect 41514 150854 42134 150938
rect 41514 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 42134 150854
rect 41514 115174 42134 150618
rect 41514 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 42134 115174
rect 41514 114854 42134 114938
rect 41514 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 42134 114854
rect 41514 79174 42134 114618
rect 41514 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 42134 79174
rect 41514 78854 42134 78938
rect 41514 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 42134 78854
rect 41514 43174 42134 78618
rect 41514 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 42134 43174
rect 41514 42854 42134 42938
rect 41514 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 42134 42854
rect 41514 7174 42134 42618
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -2266 42134 6618
rect 41514 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 42134 -2266
rect 41514 -2586 42134 -2502
rect 41514 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 42134 -2586
rect 41514 -3814 42134 -2822
rect 45234 694894 45854 708122
rect 45234 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 45854 694894
rect 45234 694574 45854 694658
rect 45234 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 45854 694574
rect 45234 658894 45854 694338
rect 45234 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 45854 658894
rect 45234 658574 45854 658658
rect 45234 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 45854 658574
rect 45234 622894 45854 658338
rect 45234 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 45854 622894
rect 45234 622574 45854 622658
rect 45234 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 45854 622574
rect 45234 586894 45854 622338
rect 45234 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 45854 586894
rect 45234 586574 45854 586658
rect 45234 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 45854 586574
rect 45234 550894 45854 586338
rect 45234 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 45854 550894
rect 45234 550574 45854 550658
rect 45234 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 45854 550574
rect 45234 514894 45854 550338
rect 45234 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 45854 514894
rect 45234 514574 45854 514658
rect 45234 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 45854 514574
rect 45234 478894 45854 514338
rect 45234 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 45854 478894
rect 45234 478574 45854 478658
rect 45234 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 45854 478574
rect 45234 442894 45854 478338
rect 48954 698614 49574 710042
rect 66954 711558 67574 711590
rect 66954 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 67574 711558
rect 66954 711238 67574 711322
rect 66954 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 67574 711238
rect 63234 709638 63854 709670
rect 63234 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 63854 709638
rect 63234 709318 63854 709402
rect 63234 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 63854 709318
rect 59514 707718 60134 707750
rect 59514 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 60134 707718
rect 59514 707398 60134 707482
rect 59514 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 60134 707398
rect 48954 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 49574 698614
rect 48954 698294 49574 698378
rect 48954 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 49574 698294
rect 48954 662614 49574 698058
rect 48954 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 49574 662614
rect 48954 662294 49574 662378
rect 48954 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 49574 662294
rect 48954 626614 49574 662058
rect 48954 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 49574 626614
rect 48954 626294 49574 626378
rect 48954 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 49574 626294
rect 48954 590614 49574 626058
rect 48954 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 49574 590614
rect 48954 590294 49574 590378
rect 48954 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 49574 590294
rect 48954 554614 49574 590058
rect 48954 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 49574 554614
rect 48954 554294 49574 554378
rect 48954 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 49574 554294
rect 48954 518614 49574 554058
rect 48954 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 49574 518614
rect 48954 518294 49574 518378
rect 48954 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 49574 518294
rect 48954 482614 49574 518058
rect 48954 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 49574 482614
rect 48954 482294 49574 482378
rect 48954 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 49574 482294
rect 48954 465308 49574 482058
rect 55794 705798 56414 705830
rect 55794 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 56414 705798
rect 55794 705478 56414 705562
rect 55794 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 56414 705478
rect 55794 669454 56414 705242
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 465308 56414 488898
rect 59514 673174 60134 707162
rect 59514 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 60134 673174
rect 59514 672854 60134 672938
rect 59514 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 60134 672854
rect 59514 637174 60134 672618
rect 59514 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 60134 637174
rect 59514 636854 60134 636938
rect 59514 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 60134 636854
rect 59514 601174 60134 636618
rect 59514 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 60134 601174
rect 59514 600854 60134 600938
rect 59514 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 60134 600854
rect 59514 565174 60134 600618
rect 59514 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 60134 565174
rect 59514 564854 60134 564938
rect 59514 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 60134 564854
rect 59514 529174 60134 564618
rect 59514 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 60134 529174
rect 59514 528854 60134 528938
rect 59514 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 60134 528854
rect 59514 493174 60134 528618
rect 59514 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 60134 493174
rect 59514 492854 60134 492938
rect 59514 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 60134 492854
rect 59514 465308 60134 492618
rect 63234 676894 63854 709082
rect 63234 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 63854 676894
rect 63234 676574 63854 676658
rect 63234 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 63854 676574
rect 63234 640894 63854 676338
rect 63234 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 63854 640894
rect 63234 640574 63854 640658
rect 63234 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 63854 640574
rect 63234 604894 63854 640338
rect 63234 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 63854 604894
rect 63234 604574 63854 604658
rect 63234 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 63854 604574
rect 63234 568894 63854 604338
rect 63234 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 63854 568894
rect 63234 568574 63854 568658
rect 63234 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 63854 568574
rect 63234 532894 63854 568338
rect 63234 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 63854 532894
rect 63234 532574 63854 532658
rect 63234 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 63854 532574
rect 63234 496894 63854 532338
rect 63234 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 63854 496894
rect 63234 496574 63854 496658
rect 63234 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 63854 496574
rect 63234 465308 63854 496338
rect 66954 680614 67574 711002
rect 84954 710598 85574 711590
rect 84954 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 85574 710598
rect 84954 710278 85574 710362
rect 84954 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 85574 710278
rect 81234 708678 81854 709670
rect 81234 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 81854 708678
rect 81234 708358 81854 708442
rect 81234 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 81854 708358
rect 77514 706758 78134 707750
rect 77514 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 78134 706758
rect 77514 706438 78134 706522
rect 77514 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 78134 706438
rect 66954 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 67574 680614
rect 66954 680294 67574 680378
rect 66954 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 67574 680294
rect 66954 644614 67574 680058
rect 66954 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 67574 644614
rect 66954 644294 67574 644378
rect 66954 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 67574 644294
rect 66954 608614 67574 644058
rect 66954 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 67574 608614
rect 66954 608294 67574 608378
rect 66954 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 67574 608294
rect 66954 572614 67574 608058
rect 66954 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 67574 572614
rect 66954 572294 67574 572378
rect 66954 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 67574 572294
rect 66954 536614 67574 572058
rect 66954 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 67574 536614
rect 66954 536294 67574 536378
rect 66954 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 67574 536294
rect 66954 500614 67574 536058
rect 66954 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 67574 500614
rect 66954 500294 67574 500378
rect 66954 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 67574 500294
rect 66954 465308 67574 500058
rect 73794 704838 74414 705830
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 579454 74414 614898
rect 73794 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 74414 579454
rect 73794 579134 74414 579218
rect 73794 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 74414 579134
rect 73794 543454 74414 578898
rect 73794 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 74414 543454
rect 73794 543134 74414 543218
rect 73794 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 74414 543134
rect 73794 507454 74414 542898
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 471454 74414 506898
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73794 465308 74414 470898
rect 77514 691174 78134 706202
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 655174 78134 690618
rect 77514 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 78134 655174
rect 77514 654854 78134 654938
rect 77514 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 78134 654854
rect 77514 619174 78134 654618
rect 77514 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 78134 619174
rect 77514 618854 78134 618938
rect 77514 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 78134 618854
rect 77514 583174 78134 618618
rect 77514 582938 77546 583174
rect 77782 582938 77866 583174
rect 78102 582938 78134 583174
rect 77514 582854 78134 582938
rect 77514 582618 77546 582854
rect 77782 582618 77866 582854
rect 78102 582618 78134 582854
rect 77514 547174 78134 582618
rect 77514 546938 77546 547174
rect 77782 546938 77866 547174
rect 78102 546938 78134 547174
rect 77514 546854 78134 546938
rect 77514 546618 77546 546854
rect 77782 546618 77866 546854
rect 78102 546618 78134 546854
rect 77514 511174 78134 546618
rect 77514 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 78134 511174
rect 77514 510854 78134 510938
rect 77514 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 78134 510854
rect 77514 475174 78134 510618
rect 77514 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 78134 475174
rect 77514 474854 78134 474938
rect 77514 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 78134 474854
rect 77514 465308 78134 474618
rect 81234 694894 81854 708122
rect 81234 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 81854 694894
rect 81234 694574 81854 694658
rect 81234 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 81854 694574
rect 81234 658894 81854 694338
rect 81234 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 81854 658894
rect 81234 658574 81854 658658
rect 81234 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 81854 658574
rect 81234 622894 81854 658338
rect 81234 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 81854 622894
rect 81234 622574 81854 622658
rect 81234 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 81854 622574
rect 81234 586894 81854 622338
rect 81234 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 81854 586894
rect 81234 586574 81854 586658
rect 81234 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 81854 586574
rect 81234 550894 81854 586338
rect 81234 550658 81266 550894
rect 81502 550658 81586 550894
rect 81822 550658 81854 550894
rect 81234 550574 81854 550658
rect 81234 550338 81266 550574
rect 81502 550338 81586 550574
rect 81822 550338 81854 550574
rect 81234 514894 81854 550338
rect 81234 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 81854 514894
rect 81234 514574 81854 514658
rect 81234 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 81854 514574
rect 81234 478894 81854 514338
rect 81234 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 81854 478894
rect 81234 478574 81854 478658
rect 81234 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 81854 478574
rect 81019 465764 81085 465765
rect 81019 465700 81020 465764
rect 81084 465700 81085 465764
rect 81019 465699 81085 465700
rect 78811 465628 78877 465629
rect 78811 465564 78812 465628
rect 78876 465564 78877 465628
rect 78811 465563 78877 465564
rect 78814 463450 78874 465563
rect 81022 463450 81082 465699
rect 81234 465308 81854 478338
rect 84954 698614 85574 710042
rect 102954 711558 103574 711590
rect 102954 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 103574 711558
rect 102954 711238 103574 711322
rect 102954 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 103574 711238
rect 99234 709638 99854 709670
rect 99234 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 99854 709638
rect 99234 709318 99854 709402
rect 99234 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 99854 709318
rect 95514 707718 96134 707750
rect 95514 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 96134 707718
rect 95514 707398 96134 707482
rect 95514 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 96134 707398
rect 84954 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 85574 698614
rect 84954 698294 85574 698378
rect 84954 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 85574 698294
rect 84954 662614 85574 698058
rect 84954 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 85574 662614
rect 84954 662294 85574 662378
rect 84954 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 85574 662294
rect 84954 626614 85574 662058
rect 84954 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 85574 626614
rect 84954 626294 85574 626378
rect 84954 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 85574 626294
rect 84954 590614 85574 626058
rect 84954 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 85574 590614
rect 84954 590294 85574 590378
rect 84954 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 85574 590294
rect 84954 554614 85574 590058
rect 84954 554378 84986 554614
rect 85222 554378 85306 554614
rect 85542 554378 85574 554614
rect 84954 554294 85574 554378
rect 84954 554058 84986 554294
rect 85222 554058 85306 554294
rect 85542 554058 85574 554294
rect 84954 518614 85574 554058
rect 84954 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 85574 518614
rect 84954 518294 85574 518378
rect 84954 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 85574 518294
rect 84954 482614 85574 518058
rect 84954 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 85574 482614
rect 84954 482294 85574 482378
rect 84954 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 85574 482294
rect 84954 465308 85574 482058
rect 91794 705798 92414 705830
rect 91794 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 92414 705798
rect 91794 705478 92414 705562
rect 91794 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 92414 705478
rect 91794 669454 92414 705242
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 91794 561454 92414 596898
rect 91794 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 92414 561454
rect 91794 561134 92414 561218
rect 91794 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 92414 561134
rect 91794 525454 92414 560898
rect 91794 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 92414 525454
rect 91794 525134 92414 525218
rect 91794 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 92414 525134
rect 91794 489454 92414 524898
rect 91794 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 92414 489454
rect 91794 489134 92414 489218
rect 91794 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 92414 489134
rect 86171 466172 86237 466173
rect 86171 466108 86172 466172
rect 86236 466108 86237 466172
rect 86171 466107 86237 466108
rect 83461 463724 83527 463725
rect 83461 463660 83462 463724
rect 83526 463660 83527 463724
rect 83461 463659 83527 463660
rect 78704 463390 78874 463450
rect 81016 463390 81082 463450
rect 78704 463202 78764 463390
rect 81016 463202 81076 463390
rect 83464 463202 83524 463659
rect 86174 463450 86234 466107
rect 88563 466036 88629 466037
rect 88563 465972 88564 466036
rect 88628 465972 88629 466036
rect 88563 465971 88629 465972
rect 88566 463450 88626 465971
rect 91794 465308 92414 488898
rect 95514 673174 96134 707162
rect 95514 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 96134 673174
rect 95514 672854 96134 672938
rect 95514 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 96134 672854
rect 95514 637174 96134 672618
rect 95514 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 96134 637174
rect 95514 636854 96134 636938
rect 95514 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 96134 636854
rect 95514 601174 96134 636618
rect 95514 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 96134 601174
rect 95514 600854 96134 600938
rect 95514 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 96134 600854
rect 95514 565174 96134 600618
rect 95514 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 96134 565174
rect 95514 564854 96134 564938
rect 95514 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 96134 564854
rect 95514 529174 96134 564618
rect 95514 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 96134 529174
rect 95514 528854 96134 528938
rect 95514 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 96134 528854
rect 95514 493174 96134 528618
rect 95514 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 96134 493174
rect 95514 492854 96134 492938
rect 95514 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 96134 492854
rect 93531 465900 93597 465901
rect 93531 465836 93532 465900
rect 93596 465836 93597 465900
rect 93531 465835 93597 465836
rect 91139 465220 91205 465221
rect 91139 465156 91140 465220
rect 91204 465156 91205 465220
rect 91139 465155 91205 465156
rect 91142 463450 91202 465155
rect 93534 463450 93594 465835
rect 95514 465308 96134 492618
rect 99234 676894 99854 709082
rect 99234 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 99854 676894
rect 99234 676574 99854 676658
rect 99234 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 99854 676574
rect 99234 640894 99854 676338
rect 99234 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 99854 640894
rect 99234 640574 99854 640658
rect 99234 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 99854 640574
rect 99234 604894 99854 640338
rect 99234 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 99854 604894
rect 99234 604574 99854 604658
rect 99234 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 99854 604574
rect 99234 568894 99854 604338
rect 99234 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 99854 568894
rect 99234 568574 99854 568658
rect 99234 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 99854 568574
rect 99234 532894 99854 568338
rect 99234 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 99854 532894
rect 99234 532574 99854 532658
rect 99234 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 99854 532574
rect 99234 496894 99854 532338
rect 99234 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 99854 496894
rect 99234 496574 99854 496658
rect 99234 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 99854 496574
rect 99234 465308 99854 496338
rect 102954 680614 103574 711002
rect 120954 710598 121574 711590
rect 120954 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 121574 710598
rect 120954 710278 121574 710362
rect 120954 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 121574 710278
rect 117234 708678 117854 709670
rect 117234 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 117854 708678
rect 117234 708358 117854 708442
rect 117234 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 117854 708358
rect 113514 706758 114134 707750
rect 113514 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 114134 706758
rect 113514 706438 114134 706522
rect 113514 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 114134 706438
rect 102954 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 103574 680614
rect 102954 680294 103574 680378
rect 102954 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 103574 680294
rect 102954 644614 103574 680058
rect 102954 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 103574 644614
rect 102954 644294 103574 644378
rect 102954 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 103574 644294
rect 102954 608614 103574 644058
rect 102954 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 103574 608614
rect 102954 608294 103574 608378
rect 102954 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 103574 608294
rect 102954 572614 103574 608058
rect 102954 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 103574 572614
rect 102954 572294 103574 572378
rect 102954 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 103574 572294
rect 102954 536614 103574 572058
rect 102954 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 103574 536614
rect 102954 536294 103574 536378
rect 102954 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 103574 536294
rect 102954 500614 103574 536058
rect 102954 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 103574 500614
rect 102954 500294 103574 500378
rect 102954 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 103574 500294
rect 102954 465308 103574 500058
rect 109794 704838 110414 705830
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 109794 543454 110414 578898
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 109794 507454 110414 542898
rect 109794 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 110414 507454
rect 109794 507134 110414 507218
rect 109794 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 110414 507134
rect 109794 471454 110414 506898
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 108435 465492 108501 465493
rect 108435 465428 108436 465492
rect 108500 465428 108501 465492
rect 108435 465427 108501 465428
rect 106227 465356 106293 465357
rect 106227 465292 106228 465356
rect 106292 465292 106293 465356
rect 106227 465291 106293 465292
rect 96107 465220 96173 465221
rect 96107 465156 96108 465220
rect 96172 465156 96173 465220
rect 96107 465155 96173 465156
rect 98499 465220 98565 465221
rect 98499 465156 98500 465220
rect 98564 465156 98565 465220
rect 98499 465155 98565 465156
rect 101259 465220 101325 465221
rect 101259 465156 101260 465220
rect 101324 465156 101325 465220
rect 101259 465155 101325 465156
rect 103651 465220 103717 465221
rect 103651 465156 103652 465220
rect 103716 465156 103717 465220
rect 103651 465155 103717 465156
rect 96110 463710 96170 465155
rect 98502 463710 98562 465155
rect 101262 463710 101322 465155
rect 96110 463650 96172 463710
rect 98502 463650 98620 463710
rect 86174 463390 86244 463450
rect 86184 463202 86244 463390
rect 88496 463390 88626 463450
rect 91080 463390 91202 463450
rect 93528 463390 93594 463450
rect 88496 463202 88556 463390
rect 91080 463202 91140 463390
rect 93528 463202 93588 463390
rect 96112 463202 96172 463650
rect 98560 463202 98620 463650
rect 101144 463650 101322 463710
rect 101144 463202 101204 463650
rect 103654 463450 103714 465155
rect 106230 463450 106290 465291
rect 103592 463390 103714 463450
rect 106176 463390 106290 463450
rect 108438 463450 108498 465427
rect 109794 465308 110414 470898
rect 113514 691174 114134 706202
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 113514 655174 114134 690618
rect 113514 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 114134 655174
rect 113514 654854 114134 654938
rect 113514 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 114134 654854
rect 113514 619174 114134 654618
rect 113514 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 114134 619174
rect 113514 618854 114134 618938
rect 113514 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 114134 618854
rect 113514 583174 114134 618618
rect 113514 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 114134 583174
rect 113514 582854 114134 582938
rect 113514 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 114134 582854
rect 113514 547174 114134 582618
rect 113514 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 114134 547174
rect 113514 546854 114134 546938
rect 113514 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 114134 546854
rect 113514 511174 114134 546618
rect 113514 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 114134 511174
rect 113514 510854 114134 510938
rect 113514 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 114134 510854
rect 113514 475174 114134 510618
rect 113514 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 114134 475174
rect 113514 474854 114134 474938
rect 113514 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 114134 474854
rect 113514 465308 114134 474618
rect 117234 694894 117854 708122
rect 117234 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 117854 694894
rect 117234 694574 117854 694658
rect 117234 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 117854 694574
rect 117234 658894 117854 694338
rect 117234 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 117854 658894
rect 117234 658574 117854 658658
rect 117234 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 117854 658574
rect 117234 622894 117854 658338
rect 117234 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 117854 622894
rect 117234 622574 117854 622658
rect 117234 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 117854 622574
rect 117234 586894 117854 622338
rect 117234 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 117854 586894
rect 117234 586574 117854 586658
rect 117234 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 117854 586574
rect 117234 550894 117854 586338
rect 117234 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 117854 550894
rect 117234 550574 117854 550658
rect 117234 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 117854 550574
rect 117234 514894 117854 550338
rect 117234 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 117854 514894
rect 117234 514574 117854 514658
rect 117234 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 117854 514574
rect 117234 478894 117854 514338
rect 117234 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 117854 478894
rect 117234 478574 117854 478658
rect 117234 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 117854 478574
rect 117234 465308 117854 478338
rect 120954 698614 121574 710042
rect 138954 711558 139574 711590
rect 138954 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 139574 711558
rect 138954 711238 139574 711322
rect 138954 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 139574 711238
rect 135234 709638 135854 709670
rect 135234 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 135854 709638
rect 135234 709318 135854 709402
rect 135234 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 135854 709318
rect 131514 707718 132134 707750
rect 131514 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 132134 707718
rect 131514 707398 132134 707482
rect 131514 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 132134 707398
rect 120954 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 121574 698614
rect 120954 698294 121574 698378
rect 120954 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 121574 698294
rect 120954 662614 121574 698058
rect 120954 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 121574 662614
rect 120954 662294 121574 662378
rect 120954 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 121574 662294
rect 120954 626614 121574 662058
rect 120954 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 121574 626614
rect 120954 626294 121574 626378
rect 120954 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 121574 626294
rect 120954 590614 121574 626058
rect 120954 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 121574 590614
rect 120954 590294 121574 590378
rect 120954 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 121574 590294
rect 120954 554614 121574 590058
rect 120954 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 121574 554614
rect 120954 554294 121574 554378
rect 120954 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 121574 554294
rect 120954 518614 121574 554058
rect 120954 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 121574 518614
rect 120954 518294 121574 518378
rect 120954 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 121574 518294
rect 120954 482614 121574 518058
rect 120954 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 121574 482614
rect 120954 482294 121574 482378
rect 120954 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 121574 482294
rect 120954 465308 121574 482058
rect 127794 705798 128414 705830
rect 127794 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 128414 705798
rect 127794 705478 128414 705562
rect 127794 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 128414 705478
rect 127794 669454 128414 705242
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 127794 561454 128414 596898
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 127794 525454 128414 560898
rect 127794 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 128414 525454
rect 127794 525134 128414 525218
rect 127794 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 128414 525134
rect 127794 489454 128414 524898
rect 127794 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 128414 489454
rect 127794 489134 128414 489218
rect 127794 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 128414 489134
rect 127794 465308 128414 488898
rect 131514 673174 132134 707162
rect 131514 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 132134 673174
rect 131514 672854 132134 672938
rect 131514 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 132134 672854
rect 131514 637174 132134 672618
rect 131514 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 132134 637174
rect 131514 636854 132134 636938
rect 131514 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 132134 636854
rect 131514 601174 132134 636618
rect 131514 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 132134 601174
rect 131514 600854 132134 600938
rect 131514 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 132134 600854
rect 131514 565174 132134 600618
rect 131514 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 132134 565174
rect 131514 564854 132134 564938
rect 131514 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 132134 564854
rect 131514 529174 132134 564618
rect 131514 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 132134 529174
rect 131514 528854 132134 528938
rect 131514 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 132134 528854
rect 131514 493174 132134 528618
rect 131514 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 132134 493174
rect 131514 492854 132134 492938
rect 131514 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 132134 492854
rect 131514 465308 132134 492618
rect 135234 676894 135854 709082
rect 135234 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 135854 676894
rect 135234 676574 135854 676658
rect 135234 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 135854 676574
rect 135234 640894 135854 676338
rect 135234 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 135854 640894
rect 135234 640574 135854 640658
rect 135234 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 135854 640574
rect 135234 604894 135854 640338
rect 135234 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 135854 604894
rect 135234 604574 135854 604658
rect 135234 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 135854 604574
rect 135234 568894 135854 604338
rect 135234 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 135854 568894
rect 135234 568574 135854 568658
rect 135234 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 135854 568574
rect 135234 532894 135854 568338
rect 135234 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 135854 532894
rect 135234 532574 135854 532658
rect 135234 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 135854 532574
rect 135234 496894 135854 532338
rect 135234 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 135854 496894
rect 135234 496574 135854 496658
rect 135234 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 135854 496574
rect 135234 465308 135854 496338
rect 138954 680614 139574 711002
rect 156954 710598 157574 711590
rect 156954 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 157574 710598
rect 156954 710278 157574 710362
rect 156954 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 157574 710278
rect 153234 708678 153854 709670
rect 153234 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 153854 708678
rect 153234 708358 153854 708442
rect 153234 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 153854 708358
rect 149514 706758 150134 707750
rect 149514 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 150134 706758
rect 149514 706438 150134 706522
rect 149514 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 150134 706438
rect 138954 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 139574 680614
rect 138954 680294 139574 680378
rect 138954 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 139574 680294
rect 138954 644614 139574 680058
rect 138954 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 139574 644614
rect 138954 644294 139574 644378
rect 138954 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 139574 644294
rect 138954 608614 139574 644058
rect 138954 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 139574 608614
rect 138954 608294 139574 608378
rect 138954 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 139574 608294
rect 138954 572614 139574 608058
rect 138954 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 139574 572614
rect 138954 572294 139574 572378
rect 138954 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 139574 572294
rect 138954 536614 139574 572058
rect 138954 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 139574 536614
rect 138954 536294 139574 536378
rect 138954 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 139574 536294
rect 138954 500614 139574 536058
rect 138954 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 139574 500614
rect 138954 500294 139574 500378
rect 138954 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 139574 500294
rect 138954 465308 139574 500058
rect 145794 704838 146414 705830
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 543454 146414 578898
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 507454 146414 542898
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 145794 471454 146414 506898
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 465308 146414 470898
rect 149514 691174 150134 706202
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 655174 150134 690618
rect 149514 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 150134 655174
rect 149514 654854 150134 654938
rect 149514 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 150134 654854
rect 149514 619174 150134 654618
rect 149514 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 150134 619174
rect 149514 618854 150134 618938
rect 149514 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 150134 618854
rect 149514 583174 150134 618618
rect 149514 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 150134 583174
rect 149514 582854 150134 582938
rect 149514 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 150134 582854
rect 149514 547174 150134 582618
rect 149514 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 150134 547174
rect 149514 546854 150134 546938
rect 149514 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 150134 546854
rect 149514 511174 150134 546618
rect 149514 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 150134 511174
rect 149514 510854 150134 510938
rect 149514 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 150134 510854
rect 149514 475174 150134 510618
rect 149514 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 150134 475174
rect 149514 474854 150134 474938
rect 149514 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 150134 474854
rect 149514 465308 150134 474618
rect 153234 694894 153854 708122
rect 153234 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 153854 694894
rect 153234 694574 153854 694658
rect 153234 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 153854 694574
rect 153234 658894 153854 694338
rect 153234 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 153854 658894
rect 153234 658574 153854 658658
rect 153234 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 153854 658574
rect 153234 622894 153854 658338
rect 153234 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 153854 622894
rect 153234 622574 153854 622658
rect 153234 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 153854 622574
rect 153234 586894 153854 622338
rect 153234 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 153854 586894
rect 153234 586574 153854 586658
rect 153234 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 153854 586574
rect 153234 550894 153854 586338
rect 153234 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 153854 550894
rect 153234 550574 153854 550658
rect 153234 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 153854 550574
rect 153234 514894 153854 550338
rect 153234 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 153854 514894
rect 153234 514574 153854 514658
rect 153234 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 153854 514574
rect 153234 478894 153854 514338
rect 153234 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 153854 478894
rect 153234 478574 153854 478658
rect 153234 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 153854 478574
rect 153234 465308 153854 478338
rect 156954 698614 157574 710042
rect 174954 711558 175574 711590
rect 174954 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 175574 711558
rect 174954 711238 175574 711322
rect 174954 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 175574 711238
rect 171234 709638 171854 709670
rect 171234 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 171854 709638
rect 171234 709318 171854 709402
rect 171234 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 171854 709318
rect 167514 707718 168134 707750
rect 167514 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 168134 707718
rect 167514 707398 168134 707482
rect 167514 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 168134 707398
rect 156954 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 157574 698614
rect 156954 698294 157574 698378
rect 156954 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 157574 698294
rect 156954 662614 157574 698058
rect 156954 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 157574 662614
rect 156954 662294 157574 662378
rect 156954 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 157574 662294
rect 156954 626614 157574 662058
rect 156954 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 157574 626614
rect 156954 626294 157574 626378
rect 156954 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 157574 626294
rect 156954 590614 157574 626058
rect 156954 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 157574 590614
rect 156954 590294 157574 590378
rect 156954 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 157574 590294
rect 156954 554614 157574 590058
rect 156954 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 157574 554614
rect 156954 554294 157574 554378
rect 156954 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 157574 554294
rect 156954 518614 157574 554058
rect 156954 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 157574 518614
rect 156954 518294 157574 518378
rect 156954 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 157574 518294
rect 156954 482614 157574 518058
rect 156954 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 157574 482614
rect 156954 482294 157574 482378
rect 156954 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 157574 482294
rect 156954 465308 157574 482058
rect 163794 705798 164414 705830
rect 163794 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 164414 705798
rect 163794 705478 164414 705562
rect 163794 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 164414 705478
rect 163794 669454 164414 705242
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 163794 561454 164414 596898
rect 163794 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 164414 561454
rect 163794 561134 164414 561218
rect 163794 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 164414 561134
rect 163794 525454 164414 560898
rect 163794 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 164414 525454
rect 163794 525134 164414 525218
rect 163794 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 164414 525134
rect 163794 489454 164414 524898
rect 163794 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 164414 489454
rect 163794 489134 164414 489218
rect 163794 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 164414 489134
rect 163794 465308 164414 488898
rect 167514 673174 168134 707162
rect 167514 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 168134 673174
rect 167514 672854 168134 672938
rect 167514 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 168134 672854
rect 167514 637174 168134 672618
rect 167514 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 168134 637174
rect 167514 636854 168134 636938
rect 167514 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 168134 636854
rect 167514 601174 168134 636618
rect 167514 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 168134 601174
rect 167514 600854 168134 600938
rect 167514 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 168134 600854
rect 167514 565174 168134 600618
rect 167514 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 168134 565174
rect 167514 564854 168134 564938
rect 167514 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 168134 564854
rect 167514 529174 168134 564618
rect 167514 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 168134 529174
rect 167514 528854 168134 528938
rect 167514 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 168134 528854
rect 167514 493174 168134 528618
rect 167514 492938 167546 493174
rect 167782 492938 167866 493174
rect 168102 492938 168134 493174
rect 167514 492854 168134 492938
rect 167514 492618 167546 492854
rect 167782 492618 167866 492854
rect 168102 492618 168134 492854
rect 167514 465308 168134 492618
rect 171234 676894 171854 709082
rect 171234 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 171854 676894
rect 171234 676574 171854 676658
rect 171234 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 171854 676574
rect 171234 640894 171854 676338
rect 171234 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 171854 640894
rect 171234 640574 171854 640658
rect 171234 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 171854 640574
rect 171234 604894 171854 640338
rect 171234 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 171854 604894
rect 171234 604574 171854 604658
rect 171234 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 171854 604574
rect 171234 568894 171854 604338
rect 171234 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 171854 568894
rect 171234 568574 171854 568658
rect 171234 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 171854 568574
rect 171234 532894 171854 568338
rect 171234 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 171854 532894
rect 171234 532574 171854 532658
rect 171234 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 171854 532574
rect 171234 496894 171854 532338
rect 171234 496658 171266 496894
rect 171502 496658 171586 496894
rect 171822 496658 171854 496894
rect 171234 496574 171854 496658
rect 171234 496338 171266 496574
rect 171502 496338 171586 496574
rect 171822 496338 171854 496574
rect 171234 465308 171854 496338
rect 174954 680614 175574 711002
rect 192954 710598 193574 711590
rect 192954 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 193574 710598
rect 192954 710278 193574 710362
rect 192954 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 193574 710278
rect 189234 708678 189854 709670
rect 189234 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 189854 708678
rect 189234 708358 189854 708442
rect 189234 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 189854 708358
rect 185514 706758 186134 707750
rect 185514 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 186134 706758
rect 185514 706438 186134 706522
rect 185514 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 186134 706438
rect 174954 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 175574 680614
rect 174954 680294 175574 680378
rect 174954 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 175574 680294
rect 174954 644614 175574 680058
rect 174954 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 175574 644614
rect 174954 644294 175574 644378
rect 174954 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 175574 644294
rect 174954 608614 175574 644058
rect 174954 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 175574 608614
rect 174954 608294 175574 608378
rect 174954 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 175574 608294
rect 174954 572614 175574 608058
rect 174954 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 175574 572614
rect 174954 572294 175574 572378
rect 174954 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 175574 572294
rect 174954 536614 175574 572058
rect 174954 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 175574 536614
rect 174954 536294 175574 536378
rect 174954 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 175574 536294
rect 174954 500614 175574 536058
rect 174954 500378 174986 500614
rect 175222 500378 175306 500614
rect 175542 500378 175574 500614
rect 174954 500294 175574 500378
rect 174954 500058 174986 500294
rect 175222 500058 175306 500294
rect 175542 500058 175574 500294
rect 174954 465308 175574 500058
rect 181794 704838 182414 705830
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 181794 471454 182414 506898
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 181794 465308 182414 470898
rect 185514 691174 186134 706202
rect 185514 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 186134 691174
rect 185514 690854 186134 690938
rect 185514 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 186134 690854
rect 185514 655174 186134 690618
rect 185514 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 186134 655174
rect 185514 654854 186134 654938
rect 185514 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 186134 654854
rect 185514 619174 186134 654618
rect 185514 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 186134 619174
rect 185514 618854 186134 618938
rect 185514 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 186134 618854
rect 185514 583174 186134 618618
rect 185514 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 186134 583174
rect 185514 582854 186134 582938
rect 185514 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 186134 582854
rect 185514 547174 186134 582618
rect 185514 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 186134 547174
rect 185514 546854 186134 546938
rect 185514 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 186134 546854
rect 185514 511174 186134 546618
rect 185514 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 186134 511174
rect 185514 510854 186134 510938
rect 185514 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 186134 510854
rect 185514 475174 186134 510618
rect 185514 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 186134 475174
rect 185514 474854 186134 474938
rect 185514 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 186134 474854
rect 185514 465308 186134 474618
rect 189234 694894 189854 708122
rect 189234 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 189854 694894
rect 189234 694574 189854 694658
rect 189234 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 189854 694574
rect 189234 658894 189854 694338
rect 189234 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 189854 658894
rect 189234 658574 189854 658658
rect 189234 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 189854 658574
rect 189234 622894 189854 658338
rect 189234 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 189854 622894
rect 189234 622574 189854 622658
rect 189234 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 189854 622574
rect 189234 586894 189854 622338
rect 189234 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 189854 586894
rect 189234 586574 189854 586658
rect 189234 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 189854 586574
rect 189234 550894 189854 586338
rect 189234 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 189854 550894
rect 189234 550574 189854 550658
rect 189234 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 189854 550574
rect 189234 514894 189854 550338
rect 189234 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 189854 514894
rect 189234 514574 189854 514658
rect 189234 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 189854 514574
rect 189234 478894 189854 514338
rect 189234 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 189854 478894
rect 189234 478574 189854 478658
rect 189234 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 189854 478574
rect 111011 465220 111077 465221
rect 111011 465156 111012 465220
rect 111076 465156 111077 465220
rect 111011 465155 111077 465156
rect 113771 465220 113837 465221
rect 113771 465156 113772 465220
rect 113836 465156 113837 465220
rect 113771 465155 113837 465156
rect 116163 465220 116229 465221
rect 116163 465156 116164 465220
rect 116228 465156 116229 465220
rect 116163 465155 116229 465156
rect 118555 465220 118621 465221
rect 118555 465156 118556 465220
rect 118620 465156 118621 465220
rect 118555 465155 118621 465156
rect 128675 465220 128741 465221
rect 128675 465156 128676 465220
rect 128740 465156 128741 465220
rect 128675 465155 128741 465156
rect 136035 465220 136101 465221
rect 136035 465156 136036 465220
rect 136100 465156 136101 465220
rect 136035 465155 136101 465156
rect 141003 465220 141069 465221
rect 141003 465156 141004 465220
rect 141068 465156 141069 465220
rect 141003 465155 141069 465156
rect 143579 465220 143645 465221
rect 143579 465156 143580 465220
rect 143644 465156 143645 465220
rect 143579 465155 143645 465156
rect 153331 465220 153397 465221
rect 153331 465156 153332 465220
rect 153396 465156 153397 465220
rect 153331 465155 153397 465156
rect 156091 465220 156157 465221
rect 156091 465156 156092 465220
rect 156156 465156 156157 465220
rect 156091 465155 156157 465156
rect 168419 465220 168485 465221
rect 168419 465156 168420 465220
rect 168484 465156 168485 465220
rect 168419 465155 168485 465156
rect 169707 465220 169773 465221
rect 169707 465156 169708 465220
rect 169772 465156 169773 465220
rect 169707 465155 169773 465156
rect 180931 465220 180997 465221
rect 180931 465156 180932 465220
rect 180996 465156 180997 465220
rect 180931 465155 180997 465156
rect 111014 463450 111074 465155
rect 113774 463450 113834 465155
rect 116166 463450 116226 465155
rect 118558 463450 118618 465155
rect 120997 463724 121063 463725
rect 120997 463660 120998 463724
rect 121062 463660 121063 463724
rect 120997 463659 121063 463660
rect 123581 463724 123647 463725
rect 123581 463660 123582 463724
rect 123646 463660 123647 463724
rect 123581 463659 123647 463660
rect 125893 463724 125959 463725
rect 125893 463660 125894 463724
rect 125958 463660 125959 463724
rect 125893 463659 125959 463660
rect 108438 463390 108548 463450
rect 103592 463202 103652 463390
rect 106176 463202 106236 463390
rect 108488 463202 108548 463390
rect 110936 463390 111074 463450
rect 113656 463390 113834 463450
rect 116104 463390 116226 463450
rect 118552 463390 118618 463450
rect 110936 463202 110996 463390
rect 113656 463202 113716 463390
rect 116104 463202 116164 463390
rect 118552 463202 118612 463390
rect 121000 463202 121060 463659
rect 123584 463202 123644 463659
rect 125896 463202 125956 463659
rect 128678 463450 128738 465155
rect 131067 463996 131133 463997
rect 131067 463932 131068 463996
rect 131132 463932 131133 463996
rect 131067 463931 131133 463932
rect 131070 463450 131130 463931
rect 133509 463724 133575 463725
rect 133509 463660 133510 463724
rect 133574 463660 133575 463724
rect 133509 463659 133575 463660
rect 128616 463390 128738 463450
rect 131064 463390 131130 463450
rect 128616 463202 128676 463390
rect 131064 463202 131124 463390
rect 133512 463202 133572 463659
rect 136038 463450 136098 465155
rect 138405 463724 138471 463725
rect 138405 463660 138406 463724
rect 138470 463660 138471 463724
rect 138405 463659 138471 463660
rect 135960 463390 136098 463450
rect 135960 463202 136020 463390
rect 138408 463202 138468 463659
rect 141006 463450 141066 465155
rect 143582 463450 143642 465155
rect 146021 463724 146087 463725
rect 146021 463660 146022 463724
rect 146086 463660 146087 463724
rect 146021 463659 146087 463660
rect 148469 463724 148535 463725
rect 148469 463660 148470 463724
rect 148534 463660 148535 463724
rect 148469 463659 148535 463660
rect 151053 463724 151119 463725
rect 151053 463660 151054 463724
rect 151118 463660 151119 463724
rect 151053 463659 151119 463660
rect 140992 463390 141066 463450
rect 143576 463390 143642 463450
rect 140992 463202 141052 463390
rect 143576 463202 143636 463390
rect 146024 463202 146084 463659
rect 148472 463202 148532 463659
rect 151056 463202 151116 463659
rect 153334 463450 153394 465155
rect 156094 463450 156154 465155
rect 153334 463390 153428 463450
rect 153368 463202 153428 463390
rect 156088 463390 156154 463450
rect 168422 463450 168482 465155
rect 169710 463450 169770 465155
rect 180934 463450 180994 465155
rect 168422 463390 168524 463450
rect 156088 463202 156148 463390
rect 168464 463202 168524 463390
rect 169688 463390 169770 463450
rect 180840 463390 180994 463450
rect 169688 463202 169748 463390
rect 180840 463202 180900 463390
rect 50272 453454 50620 453486
rect 50272 453218 50328 453454
rect 50564 453218 50620 453454
rect 50272 453134 50620 453218
rect 50272 452898 50328 453134
rect 50564 452898 50620 453134
rect 50272 452866 50620 452898
rect 186000 453454 186348 453486
rect 186000 453218 186056 453454
rect 186292 453218 186348 453454
rect 186000 453134 186348 453218
rect 186000 452898 186056 453134
rect 186292 452898 186348 453134
rect 186000 452866 186348 452898
rect 45234 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 45854 442894
rect 45234 442574 45854 442658
rect 45234 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 45854 442574
rect 45234 406894 45854 442338
rect 189234 442894 189854 478338
rect 189234 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 189854 442894
rect 189234 442574 189854 442658
rect 189234 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 189854 442574
rect 50952 435454 51300 435486
rect 50952 435218 51008 435454
rect 51244 435218 51300 435454
rect 50952 435134 51300 435218
rect 50952 434898 51008 435134
rect 51244 434898 51300 435134
rect 50952 434866 51300 434898
rect 185320 435454 185668 435486
rect 185320 435218 185376 435454
rect 185612 435218 185668 435454
rect 185320 435134 185668 435218
rect 185320 434898 185376 435134
rect 185612 434898 185668 435134
rect 185320 434866 185668 434898
rect 50272 417454 50620 417486
rect 50272 417218 50328 417454
rect 50564 417218 50620 417454
rect 50272 417134 50620 417218
rect 50272 416898 50328 417134
rect 50564 416898 50620 417134
rect 50272 416866 50620 416898
rect 186000 417454 186348 417486
rect 186000 417218 186056 417454
rect 186292 417218 186348 417454
rect 186000 417134 186348 417218
rect 186000 416898 186056 417134
rect 186292 416898 186348 417134
rect 186000 416866 186348 416898
rect 45234 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 45854 406894
rect 45234 406574 45854 406658
rect 45234 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 45854 406574
rect 45234 370894 45854 406338
rect 189234 406894 189854 442338
rect 189234 406658 189266 406894
rect 189502 406658 189586 406894
rect 189822 406658 189854 406894
rect 189234 406574 189854 406658
rect 189234 406338 189266 406574
rect 189502 406338 189586 406574
rect 189822 406338 189854 406574
rect 50952 399454 51300 399486
rect 50952 399218 51008 399454
rect 51244 399218 51300 399454
rect 50952 399134 51300 399218
rect 50952 398898 51008 399134
rect 51244 398898 51300 399134
rect 50952 398866 51300 398898
rect 185320 399454 185668 399486
rect 185320 399218 185376 399454
rect 185612 399218 185668 399454
rect 185320 399134 185668 399218
rect 185320 398898 185376 399134
rect 185612 398898 185668 399134
rect 185320 398866 185668 398898
rect 50272 381454 50620 381486
rect 50272 381218 50328 381454
rect 50564 381218 50620 381454
rect 50272 381134 50620 381218
rect 50272 380898 50328 381134
rect 50564 380898 50620 381134
rect 50272 380866 50620 380898
rect 186000 381454 186348 381486
rect 186000 381218 186056 381454
rect 186292 381218 186348 381454
rect 186000 381134 186348 381218
rect 186000 380898 186056 381134
rect 186292 380898 186348 381134
rect 186000 380866 186348 380898
rect 66056 379810 66116 380106
rect 67144 379810 67204 380106
rect 68232 379810 68292 380106
rect 69592 379810 69652 380106
rect 70544 379810 70604 380106
rect 66056 379750 66178 379810
rect 67144 379750 67282 379810
rect 68232 379750 68386 379810
rect 69592 379750 69674 379810
rect 45234 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 45854 370894
rect 45234 370574 45854 370658
rect 45234 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 45854 370574
rect 45234 334894 45854 370338
rect 45234 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 45854 334894
rect 45234 334574 45854 334658
rect 45234 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 45854 334574
rect 45234 298894 45854 334338
rect 45234 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 45854 298894
rect 45234 298574 45854 298658
rect 45234 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 45854 298574
rect 45234 262894 45854 298338
rect 48954 374614 49574 378000
rect 48954 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 49574 374614
rect 48954 374294 49574 374378
rect 48954 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 49574 374294
rect 48954 338614 49574 374058
rect 48954 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 49574 338614
rect 48954 338294 49574 338378
rect 48954 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 49574 338294
rect 48954 302614 49574 338058
rect 48954 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 49574 302614
rect 48954 302294 49574 302378
rect 48954 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 49574 302294
rect 48954 285308 49574 302058
rect 55794 345454 56414 378000
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 285308 56414 308898
rect 59514 349174 60134 378000
rect 59514 348938 59546 349174
rect 59782 348938 59866 349174
rect 60102 348938 60134 349174
rect 59514 348854 60134 348938
rect 59514 348618 59546 348854
rect 59782 348618 59866 348854
rect 60102 348618 60134 348854
rect 59514 313174 60134 348618
rect 59514 312938 59546 313174
rect 59782 312938 59866 313174
rect 60102 312938 60134 313174
rect 59514 312854 60134 312938
rect 59514 312618 59546 312854
rect 59782 312618 59866 312854
rect 60102 312618 60134 312854
rect 59514 285308 60134 312618
rect 63234 352894 63854 378000
rect 66118 377093 66178 379750
rect 67222 378181 67282 379750
rect 67219 378180 67285 378181
rect 67219 378116 67220 378180
rect 67284 378116 67285 378180
rect 67219 378115 67285 378116
rect 66115 377092 66181 377093
rect 66115 377028 66116 377092
rect 66180 377028 66181 377092
rect 66115 377027 66181 377028
rect 63234 352658 63266 352894
rect 63502 352658 63586 352894
rect 63822 352658 63854 352894
rect 63234 352574 63854 352658
rect 63234 352338 63266 352574
rect 63502 352338 63586 352574
rect 63822 352338 63854 352574
rect 63234 316894 63854 352338
rect 63234 316658 63266 316894
rect 63502 316658 63586 316894
rect 63822 316658 63854 316894
rect 63234 316574 63854 316658
rect 63234 316338 63266 316574
rect 63502 316338 63586 316574
rect 63822 316338 63854 316574
rect 63234 285308 63854 316338
rect 66954 356614 67574 378000
rect 68326 377093 68386 379750
rect 69614 377093 69674 379750
rect 70534 379750 70604 379810
rect 71768 379810 71828 380106
rect 73128 379810 73188 380106
rect 74216 379810 74276 380106
rect 71768 379750 71882 379810
rect 70534 377093 70594 379750
rect 71822 377093 71882 379750
rect 73110 379750 73188 379810
rect 74214 379750 74276 379810
rect 75440 379810 75500 380106
rect 76528 379810 76588 380106
rect 77616 379810 77676 380106
rect 78296 379810 78356 380106
rect 75440 379750 75562 379810
rect 76528 379750 76666 379810
rect 77616 379750 77770 379810
rect 73110 378045 73170 379750
rect 74214 378181 74274 379750
rect 74211 378180 74277 378181
rect 74211 378116 74212 378180
rect 74276 378116 74277 378180
rect 74211 378115 74277 378116
rect 73107 378044 73173 378045
rect 73107 377980 73108 378044
rect 73172 377980 73173 378044
rect 73107 377979 73173 377980
rect 68323 377092 68389 377093
rect 68323 377028 68324 377092
rect 68388 377028 68389 377092
rect 68323 377027 68389 377028
rect 69611 377092 69677 377093
rect 69611 377028 69612 377092
rect 69676 377028 69677 377092
rect 69611 377027 69677 377028
rect 70531 377092 70597 377093
rect 70531 377028 70532 377092
rect 70596 377028 70597 377092
rect 70531 377027 70597 377028
rect 71819 377092 71885 377093
rect 71819 377028 71820 377092
rect 71884 377028 71885 377092
rect 71819 377027 71885 377028
rect 66954 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 67574 356614
rect 66954 356294 67574 356378
rect 66954 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 67574 356294
rect 66954 320614 67574 356058
rect 66954 320378 66986 320614
rect 67222 320378 67306 320614
rect 67542 320378 67574 320614
rect 66954 320294 67574 320378
rect 66954 320058 66986 320294
rect 67222 320058 67306 320294
rect 67542 320058 67574 320294
rect 66954 285308 67574 320058
rect 73794 363454 74414 378000
rect 75502 377093 75562 379750
rect 76606 377093 76666 379750
rect 77710 378181 77770 379750
rect 78262 379750 78356 379810
rect 78704 379810 78764 380106
rect 80064 379810 80124 380106
rect 80744 379810 80804 380106
rect 81288 379810 81348 380106
rect 78704 379750 78874 379810
rect 80064 379750 80162 379810
rect 80744 379750 80898 379810
rect 77707 378180 77773 378181
rect 77707 378116 77708 378180
rect 77772 378116 77773 378180
rect 77707 378115 77773 378116
rect 75499 377092 75565 377093
rect 75499 377028 75500 377092
rect 75564 377028 75565 377092
rect 75499 377027 75565 377028
rect 76603 377092 76669 377093
rect 76603 377028 76604 377092
rect 76668 377028 76669 377092
rect 76603 377027 76669 377028
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 73794 327454 74414 362898
rect 73794 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 74414 327454
rect 73794 327134 74414 327218
rect 73794 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 74414 327134
rect 73794 291454 74414 326898
rect 73794 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 74414 291454
rect 73794 291134 74414 291218
rect 73794 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 74414 291134
rect 73794 285308 74414 290898
rect 77514 367174 78134 378000
rect 78262 377093 78322 379750
rect 78814 377093 78874 379750
rect 80102 377093 80162 379750
rect 78259 377092 78325 377093
rect 78259 377028 78260 377092
rect 78324 377028 78325 377092
rect 78259 377027 78325 377028
rect 78811 377092 78877 377093
rect 78811 377028 78812 377092
rect 78876 377028 78877 377092
rect 78811 377027 78877 377028
rect 80099 377092 80165 377093
rect 80099 377028 80100 377092
rect 80164 377028 80165 377092
rect 80099 377027 80165 377028
rect 80838 376957 80898 379750
rect 81206 379750 81348 379810
rect 82376 379810 82436 380106
rect 83464 379810 83524 380106
rect 83600 379810 83660 380106
rect 82376 379750 82554 379810
rect 81206 378181 81266 379750
rect 81203 378180 81269 378181
rect 81203 378116 81204 378180
rect 81268 378116 81269 378180
rect 81203 378115 81269 378116
rect 80835 376956 80901 376957
rect 80835 376892 80836 376956
rect 80900 376892 80901 376956
rect 80835 376891 80901 376892
rect 77514 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 78134 367174
rect 77514 366854 78134 366938
rect 77514 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 78134 366854
rect 77514 331174 78134 366618
rect 77514 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 78134 331174
rect 77514 330854 78134 330938
rect 77514 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 78134 330854
rect 77514 295174 78134 330618
rect 77514 294938 77546 295174
rect 77782 294938 77866 295174
rect 78102 294938 78134 295174
rect 77514 294854 78134 294938
rect 77514 294618 77546 294854
rect 77782 294618 77866 294854
rect 78102 294618 78134 294854
rect 77514 285308 78134 294618
rect 81234 370894 81854 378000
rect 82494 377093 82554 379750
rect 83414 379750 83524 379810
rect 83598 379750 83660 379810
rect 82491 377092 82557 377093
rect 82491 377028 82492 377092
rect 82556 377028 82557 377092
rect 82491 377027 82557 377028
rect 83414 376957 83474 379750
rect 83598 377093 83658 379750
rect 84552 379538 84612 380106
rect 85912 379810 85972 380106
rect 84518 379478 84612 379538
rect 85806 379750 85972 379810
rect 84518 377093 84578 379478
rect 83595 377092 83661 377093
rect 83595 377028 83596 377092
rect 83660 377028 83661 377092
rect 83595 377027 83661 377028
rect 84515 377092 84581 377093
rect 84515 377028 84516 377092
rect 84580 377028 84581 377092
rect 84515 377027 84581 377028
rect 83411 376956 83477 376957
rect 83411 376892 83412 376956
rect 83476 376892 83477 376956
rect 83411 376891 83477 376892
rect 81234 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 81854 370894
rect 81234 370574 81854 370658
rect 81234 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 81854 370574
rect 81234 334894 81854 370338
rect 81234 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 81854 334894
rect 81234 334574 81854 334658
rect 81234 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 81854 334574
rect 81234 298894 81854 334338
rect 81234 298658 81266 298894
rect 81502 298658 81586 298894
rect 81822 298658 81854 298894
rect 81234 298574 81854 298658
rect 81234 298338 81266 298574
rect 81502 298338 81586 298574
rect 81822 298338 81854 298574
rect 78811 286108 78877 286109
rect 78811 286044 78812 286108
rect 78876 286044 78877 286108
rect 78811 286043 78877 286044
rect 78814 283930 78874 286043
rect 81019 285836 81085 285837
rect 81019 285772 81020 285836
rect 81084 285772 81085 285836
rect 81019 285771 81085 285772
rect 81022 283930 81082 285771
rect 81234 285308 81854 298338
rect 84954 374614 85574 378000
rect 85806 376957 85866 379750
rect 86048 379538 86108 380106
rect 87000 379810 87060 380106
rect 88088 379810 88148 380106
rect 87000 379750 87154 379810
rect 85990 379478 86108 379538
rect 85990 377093 86050 379478
rect 85987 377092 86053 377093
rect 85987 377028 85988 377092
rect 86052 377028 86053 377092
rect 85987 377027 86053 377028
rect 87094 376957 87154 379750
rect 88014 379750 88148 379810
rect 88496 379810 88556 380106
rect 88496 379750 88626 379810
rect 88014 377093 88074 379750
rect 88011 377092 88077 377093
rect 88011 377028 88012 377092
rect 88076 377028 88077 377092
rect 88011 377027 88077 377028
rect 88566 376957 88626 379750
rect 89448 379538 89508 380106
rect 90672 379810 90732 380106
rect 90672 379750 90834 379810
rect 89448 379478 89546 379538
rect 89486 377093 89546 379478
rect 90774 377093 90834 379750
rect 91080 379538 91140 380106
rect 91760 379810 91820 380106
rect 91760 379750 91938 379810
rect 91080 379478 91202 379538
rect 91142 377093 91202 379478
rect 91878 378181 91938 379750
rect 92848 379538 92908 380106
rect 92798 379478 92908 379538
rect 93528 379538 93588 380106
rect 93936 379541 93996 380106
rect 93933 379540 93999 379541
rect 93528 379478 93594 379538
rect 91875 378180 91941 378181
rect 91875 378116 91876 378180
rect 91940 378116 91941 378180
rect 91875 378115 91941 378116
rect 92798 378045 92858 379478
rect 92795 378044 92861 378045
rect 89483 377092 89549 377093
rect 89483 377028 89484 377092
rect 89548 377028 89549 377092
rect 89483 377027 89549 377028
rect 90771 377092 90837 377093
rect 90771 377028 90772 377092
rect 90836 377028 90837 377092
rect 90771 377027 90837 377028
rect 91139 377092 91205 377093
rect 91139 377028 91140 377092
rect 91204 377028 91205 377092
rect 91139 377027 91205 377028
rect 85803 376956 85869 376957
rect 85803 376892 85804 376956
rect 85868 376892 85869 376956
rect 85803 376891 85869 376892
rect 87091 376956 87157 376957
rect 87091 376892 87092 376956
rect 87156 376892 87157 376956
rect 87091 376891 87157 376892
rect 88563 376956 88629 376957
rect 88563 376892 88564 376956
rect 88628 376892 88629 376956
rect 88563 376891 88629 376892
rect 84954 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 85574 374614
rect 84954 374294 85574 374378
rect 84954 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 85574 374294
rect 84954 338614 85574 374058
rect 84954 338378 84986 338614
rect 85222 338378 85306 338614
rect 85542 338378 85574 338614
rect 84954 338294 85574 338378
rect 84954 338058 84986 338294
rect 85222 338058 85306 338294
rect 85542 338058 85574 338294
rect 84954 302614 85574 338058
rect 84954 302378 84986 302614
rect 85222 302378 85306 302614
rect 85542 302378 85574 302614
rect 84954 302294 85574 302378
rect 84954 302058 84986 302294
rect 85222 302058 85306 302294
rect 85542 302058 85574 302294
rect 83411 285700 83477 285701
rect 83411 285636 83412 285700
rect 83476 285636 83477 285700
rect 83411 285635 83477 285636
rect 78704 283870 78874 283930
rect 81016 283870 81082 283930
rect 83414 283930 83474 285635
rect 84954 285308 85574 302058
rect 91794 345454 92414 378000
rect 92795 377980 92796 378044
rect 92860 377980 92861 378044
rect 92795 377979 92861 377980
rect 93534 377093 93594 379478
rect 93933 379476 93934 379540
rect 93998 379476 93999 379540
rect 95296 379530 95356 380106
rect 95976 379530 96036 380106
rect 96384 379541 96444 380106
rect 97608 379541 97668 380106
rect 93933 379475 93999 379476
rect 95190 379470 95356 379530
rect 95926 379470 96036 379530
rect 96381 379540 96447 379541
rect 96381 379476 96382 379540
rect 96446 379476 96447 379540
rect 96381 379475 96447 379476
rect 97605 379540 97671 379541
rect 97605 379476 97606 379540
rect 97670 379476 97671 379540
rect 97605 379475 97671 379476
rect 98288 379530 98348 380106
rect 98696 379541 98756 380106
rect 98693 379540 98759 379541
rect 98288 379470 98378 379530
rect 98693 379476 98694 379540
rect 98758 379476 98759 379540
rect 98693 379475 98759 379476
rect 99784 379530 99844 380106
rect 101008 379530 101068 380106
rect 101144 379810 101204 380106
rect 101144 379750 101322 379810
rect 99784 379470 99850 379530
rect 101008 379470 101138 379530
rect 95190 378045 95250 379470
rect 95926 378181 95986 379470
rect 95923 378180 95989 378181
rect 95923 378116 95924 378180
rect 95988 378116 95989 378180
rect 95923 378115 95989 378116
rect 95187 378044 95253 378045
rect 95187 377980 95188 378044
rect 95252 377980 95253 378044
rect 95187 377979 95253 377980
rect 93531 377092 93597 377093
rect 93531 377028 93532 377092
rect 93596 377028 93597 377092
rect 93531 377027 93597 377028
rect 91794 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 92414 345454
rect 91794 345134 92414 345218
rect 91794 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 92414 345134
rect 91794 309454 92414 344898
rect 91794 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 92414 309454
rect 91794 309134 92414 309218
rect 91794 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 92414 309134
rect 86171 285700 86237 285701
rect 86171 285636 86172 285700
rect 86236 285636 86237 285700
rect 86171 285635 86237 285636
rect 88563 285700 88629 285701
rect 88563 285636 88564 285700
rect 88628 285636 88629 285700
rect 88563 285635 88629 285636
rect 91139 285700 91205 285701
rect 91139 285636 91140 285700
rect 91204 285636 91205 285700
rect 91139 285635 91205 285636
rect 86174 283930 86234 285635
rect 88566 283930 88626 285635
rect 91142 283930 91202 285635
rect 91794 285308 92414 308898
rect 95514 349174 96134 378000
rect 98318 377093 98378 379470
rect 99790 378181 99850 379470
rect 99787 378180 99853 378181
rect 99787 378116 99788 378180
rect 99852 378116 99853 378180
rect 99787 378115 99853 378116
rect 98315 377092 98381 377093
rect 98315 377028 98316 377092
rect 98380 377028 98381 377092
rect 98315 377027 98381 377028
rect 95514 348938 95546 349174
rect 95782 348938 95866 349174
rect 96102 348938 96134 349174
rect 95514 348854 96134 348938
rect 95514 348618 95546 348854
rect 95782 348618 95866 348854
rect 96102 348618 96134 348854
rect 95514 313174 96134 348618
rect 95514 312938 95546 313174
rect 95782 312938 95866 313174
rect 96102 312938 96134 313174
rect 95514 312854 96134 312938
rect 95514 312618 95546 312854
rect 95782 312618 95866 312854
rect 96102 312618 96134 312854
rect 93531 285700 93597 285701
rect 93531 285636 93532 285700
rect 93596 285636 93597 285700
rect 93531 285635 93597 285636
rect 93534 283930 93594 285635
rect 95514 285308 96134 312618
rect 99234 352894 99854 378000
rect 101078 377093 101138 379470
rect 101262 378045 101322 379750
rect 102232 379541 102292 380106
rect 102229 379540 102295 379541
rect 102229 379476 102230 379540
rect 102294 379476 102295 379540
rect 103320 379530 103380 380106
rect 102229 379475 102295 379476
rect 103286 379470 103380 379530
rect 103592 379530 103652 380106
rect 104408 379530 104468 380106
rect 103592 379470 103714 379530
rect 103286 378181 103346 379470
rect 103654 378181 103714 379470
rect 104390 379470 104468 379530
rect 105768 379530 105828 380106
rect 106040 379530 106100 380106
rect 106992 379530 107052 380106
rect 108080 379810 108140 380106
rect 105768 379470 105922 379530
rect 106040 379470 106106 379530
rect 103283 378180 103349 378181
rect 103283 378116 103284 378180
rect 103348 378116 103349 378180
rect 103283 378115 103349 378116
rect 103651 378180 103717 378181
rect 103651 378116 103652 378180
rect 103716 378116 103717 378180
rect 103651 378115 103717 378116
rect 101259 378044 101325 378045
rect 101259 377980 101260 378044
rect 101324 377980 101325 378044
rect 101259 377979 101325 377980
rect 101075 377092 101141 377093
rect 101075 377028 101076 377092
rect 101140 377028 101141 377092
rect 101075 377027 101141 377028
rect 99234 352658 99266 352894
rect 99502 352658 99586 352894
rect 99822 352658 99854 352894
rect 99234 352574 99854 352658
rect 99234 352338 99266 352574
rect 99502 352338 99586 352574
rect 99822 352338 99854 352574
rect 99234 316894 99854 352338
rect 99234 316658 99266 316894
rect 99502 316658 99586 316894
rect 99822 316658 99854 316894
rect 99234 316574 99854 316658
rect 99234 316338 99266 316574
rect 99502 316338 99586 316574
rect 99822 316338 99854 316574
rect 96291 285700 96357 285701
rect 96291 285636 96292 285700
rect 96356 285636 96357 285700
rect 96291 285635 96357 285636
rect 96294 283930 96354 285635
rect 99234 285308 99854 316338
rect 102954 356614 103574 378000
rect 104390 377909 104450 379470
rect 105862 378045 105922 379470
rect 105859 378044 105925 378045
rect 105859 377980 105860 378044
rect 105924 377980 105925 378044
rect 105859 377979 105925 377980
rect 104387 377908 104453 377909
rect 104387 377844 104388 377908
rect 104452 377844 104453 377908
rect 104387 377843 104453 377844
rect 106046 377093 106106 379470
rect 106966 379470 107052 379530
rect 108070 379750 108140 379810
rect 106966 378045 107026 379470
rect 108070 379405 108130 379750
rect 108488 379530 108548 380106
rect 108438 379470 108548 379530
rect 109168 379530 109228 380106
rect 110936 379530 110996 380106
rect 113520 379810 113580 380106
rect 115968 379810 116028 380106
rect 118280 379810 118340 380106
rect 121000 379810 121060 380106
rect 113520 379750 113650 379810
rect 115968 379750 116042 379810
rect 118280 379750 118434 379810
rect 109168 379470 109234 379530
rect 110936 379470 111074 379530
rect 108067 379404 108133 379405
rect 108067 379340 108068 379404
rect 108132 379340 108133 379404
rect 108067 379339 108133 379340
rect 106963 378044 107029 378045
rect 106963 377980 106964 378044
rect 107028 377980 107029 378044
rect 106963 377979 107029 377980
rect 108438 377093 108498 379470
rect 109174 378045 109234 379470
rect 109171 378044 109237 378045
rect 109171 377980 109172 378044
rect 109236 377980 109237 378044
rect 109171 377979 109237 377980
rect 106043 377092 106109 377093
rect 106043 377028 106044 377092
rect 106108 377028 106109 377092
rect 106043 377027 106109 377028
rect 108435 377092 108501 377093
rect 108435 377028 108436 377092
rect 108500 377028 108501 377092
rect 108435 377027 108501 377028
rect 102954 356378 102986 356614
rect 103222 356378 103306 356614
rect 103542 356378 103574 356614
rect 102954 356294 103574 356378
rect 102954 356058 102986 356294
rect 103222 356058 103306 356294
rect 103542 356058 103574 356294
rect 102954 320614 103574 356058
rect 102954 320378 102986 320614
rect 103222 320378 103306 320614
rect 103542 320378 103574 320614
rect 102954 320294 103574 320378
rect 102954 320058 102986 320294
rect 103222 320058 103306 320294
rect 103542 320058 103574 320294
rect 102954 285308 103574 320058
rect 109794 363454 110414 378000
rect 111014 377093 111074 379470
rect 113590 378181 113650 379750
rect 113587 378180 113653 378181
rect 113587 378116 113588 378180
rect 113652 378116 113653 378180
rect 113587 378115 113653 378116
rect 111011 377092 111077 377093
rect 111011 377028 111012 377092
rect 111076 377028 111077 377092
rect 111011 377027 111077 377028
rect 109794 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 110414 363454
rect 109794 363134 110414 363218
rect 109794 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 110414 363134
rect 109794 327454 110414 362898
rect 109794 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 110414 327454
rect 109794 327134 110414 327218
rect 109794 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 110414 327134
rect 109794 291454 110414 326898
rect 109794 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 110414 291454
rect 109794 291134 110414 291218
rect 109794 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 110414 291134
rect 106227 285972 106293 285973
rect 106227 285908 106228 285972
rect 106292 285908 106293 285972
rect 106227 285907 106293 285908
rect 108435 285972 108501 285973
rect 108435 285908 108436 285972
rect 108500 285908 108501 285972
rect 108435 285907 108501 285908
rect 103835 285700 103901 285701
rect 103835 285636 103836 285700
rect 103900 285636 103901 285700
rect 103835 285635 103901 285636
rect 98499 284884 98565 284885
rect 98499 284820 98500 284884
rect 98564 284820 98565 284884
rect 98499 284819 98565 284820
rect 83414 283870 83524 283930
rect 86174 283870 86244 283930
rect 78704 283220 78764 283870
rect 81016 283220 81076 283870
rect 83464 283220 83524 283870
rect 86184 283220 86244 283870
rect 88496 283870 88626 283930
rect 91080 283870 91202 283930
rect 93528 283870 93594 283930
rect 96112 283870 96354 283930
rect 98502 283930 98562 284819
rect 101259 284748 101325 284749
rect 101259 284684 101260 284748
rect 101324 284684 101325 284748
rect 101259 284683 101325 284684
rect 101262 283930 101322 284683
rect 103838 283930 103898 285635
rect 106230 283930 106290 285907
rect 98502 283870 98620 283930
rect 88496 283220 88556 283870
rect 91080 283220 91140 283870
rect 93528 283220 93588 283870
rect 96112 283220 96172 283870
rect 98560 283220 98620 283870
rect 101144 283870 101322 283930
rect 103592 283870 103898 283930
rect 106176 283870 106290 283930
rect 108438 283930 108498 285907
rect 109794 285308 110414 290898
rect 113514 367174 114134 378000
rect 115982 377093 116042 379750
rect 115979 377092 116045 377093
rect 115979 377028 115980 377092
rect 116044 377028 116045 377092
rect 115979 377027 116045 377028
rect 113514 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 114134 367174
rect 113514 366854 114134 366938
rect 113514 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 114134 366854
rect 113514 331174 114134 366618
rect 113514 330938 113546 331174
rect 113782 330938 113866 331174
rect 114102 330938 114134 331174
rect 113514 330854 114134 330938
rect 113514 330618 113546 330854
rect 113782 330618 113866 330854
rect 114102 330618 114134 330854
rect 113514 295174 114134 330618
rect 113514 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 114134 295174
rect 113514 294854 114134 294938
rect 113514 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 114134 294854
rect 113514 285308 114134 294618
rect 117234 370894 117854 378000
rect 118374 377093 118434 379750
rect 120950 379750 121060 379810
rect 120950 378181 121010 379750
rect 123448 379677 123508 380106
rect 125896 379810 125956 380106
rect 128480 379810 128540 380106
rect 125896 379750 125978 379810
rect 128480 379750 128554 379810
rect 123445 379676 123511 379677
rect 123445 379612 123446 379676
rect 123510 379612 123511 379676
rect 123445 379611 123511 379612
rect 125918 379541 125978 379750
rect 128494 379541 128554 379750
rect 130928 379677 130988 380106
rect 133512 379677 133572 380106
rect 135960 379810 136020 380106
rect 138544 379810 138604 380106
rect 140992 379810 141052 380106
rect 143440 379810 143500 380106
rect 135960 379750 136098 379810
rect 138544 379750 138674 379810
rect 140992 379750 141066 379810
rect 130925 379676 130991 379677
rect 130925 379612 130926 379676
rect 130990 379612 130991 379676
rect 130925 379611 130991 379612
rect 133509 379676 133575 379677
rect 133509 379612 133510 379676
rect 133574 379612 133575 379676
rect 133509 379611 133575 379612
rect 125915 379540 125981 379541
rect 125915 379476 125916 379540
rect 125980 379476 125981 379540
rect 125915 379475 125981 379476
rect 128491 379540 128557 379541
rect 128491 379476 128492 379540
rect 128556 379476 128557 379540
rect 128491 379475 128557 379476
rect 120947 378180 121013 378181
rect 120947 378116 120948 378180
rect 121012 378116 121013 378180
rect 120947 378115 121013 378116
rect 136038 378045 136098 379750
rect 138614 378045 138674 379750
rect 141006 378045 141066 379750
rect 143398 379750 143500 379810
rect 143398 378045 143458 379750
rect 145888 379677 145948 380106
rect 148472 379677 148532 380106
rect 150920 379810 150980 380106
rect 153368 379810 153428 380106
rect 150920 379750 151002 379810
rect 145885 379676 145951 379677
rect 145885 379612 145886 379676
rect 145950 379612 145951 379676
rect 145885 379611 145951 379612
rect 148469 379676 148535 379677
rect 148469 379612 148470 379676
rect 148534 379612 148535 379676
rect 148469 379611 148535 379612
rect 150942 379269 151002 379750
rect 153334 379750 153428 379810
rect 150939 379268 151005 379269
rect 150939 379204 150940 379268
rect 151004 379204 151005 379268
rect 150939 379203 151005 379204
rect 153334 378181 153394 379750
rect 155952 379677 156012 380106
rect 173224 379810 173284 380106
rect 173206 379750 173284 379810
rect 173360 379810 173420 380106
rect 173360 379750 173450 379810
rect 155949 379676 156015 379677
rect 155949 379612 155950 379676
rect 156014 379612 156015 379676
rect 155949 379611 156015 379612
rect 153331 378180 153397 378181
rect 153331 378116 153332 378180
rect 153396 378116 153397 378180
rect 153331 378115 153397 378116
rect 136035 378044 136101 378045
rect 118371 377092 118437 377093
rect 118371 377028 118372 377092
rect 118436 377028 118437 377092
rect 118371 377027 118437 377028
rect 117234 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 117854 370894
rect 117234 370574 117854 370658
rect 117234 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 117854 370574
rect 117234 334894 117854 370338
rect 117234 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 117854 334894
rect 117234 334574 117854 334658
rect 117234 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 117854 334574
rect 117234 298894 117854 334338
rect 117234 298658 117266 298894
rect 117502 298658 117586 298894
rect 117822 298658 117854 298894
rect 117234 298574 117854 298658
rect 117234 298338 117266 298574
rect 117502 298338 117586 298574
rect 117822 298338 117854 298574
rect 114323 285700 114389 285701
rect 114323 285636 114324 285700
rect 114388 285636 114389 285700
rect 114323 285635 114389 285636
rect 111011 285020 111077 285021
rect 111011 284956 111012 285020
rect 111076 284956 111077 285020
rect 111011 284955 111077 284956
rect 111014 283930 111074 284955
rect 114326 283930 114386 285635
rect 117234 285308 117854 298338
rect 120954 374614 121574 378000
rect 120954 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 121574 374614
rect 120954 374294 121574 374378
rect 120954 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 121574 374294
rect 120954 338614 121574 374058
rect 120954 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 121574 338614
rect 120954 338294 121574 338378
rect 120954 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 121574 338294
rect 120954 302614 121574 338058
rect 120954 302378 120986 302614
rect 121222 302378 121306 302614
rect 121542 302378 121574 302614
rect 120954 302294 121574 302378
rect 120954 302058 120986 302294
rect 121222 302058 121306 302294
rect 121542 302058 121574 302294
rect 120763 285972 120829 285973
rect 120763 285908 120764 285972
rect 120828 285908 120829 285972
rect 120763 285907 120829 285908
rect 118555 285700 118621 285701
rect 118555 285636 118556 285700
rect 118620 285636 118621 285700
rect 118555 285635 118621 285636
rect 116163 285020 116229 285021
rect 116163 284956 116164 285020
rect 116228 284956 116229 285020
rect 116163 284955 116229 284956
rect 116166 283930 116226 284955
rect 118558 283930 118618 285635
rect 108438 283870 108548 283930
rect 101144 283220 101204 283870
rect 103592 283220 103652 283870
rect 106176 283220 106236 283870
rect 108488 283220 108548 283870
rect 110936 283870 111074 283930
rect 113656 283870 114386 283930
rect 116104 283870 116226 283930
rect 118552 283870 118618 283930
rect 120766 283930 120826 285907
rect 120954 285308 121574 302058
rect 127794 345454 128414 378000
rect 127794 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 128414 345454
rect 127794 345134 128414 345218
rect 127794 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 128414 345134
rect 127794 309454 128414 344898
rect 127794 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 128414 309454
rect 127794 309134 128414 309218
rect 127794 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 128414 309134
rect 123523 285700 123589 285701
rect 123523 285636 123524 285700
rect 123588 285636 123589 285700
rect 123523 285635 123589 285636
rect 125915 285700 125981 285701
rect 125915 285636 125916 285700
rect 125980 285636 125981 285700
rect 125915 285635 125981 285636
rect 123526 283930 123586 285635
rect 125918 283930 125978 285635
rect 127794 285308 128414 308898
rect 131514 349174 132134 378000
rect 131514 348938 131546 349174
rect 131782 348938 131866 349174
rect 132102 348938 132134 349174
rect 131514 348854 132134 348938
rect 131514 348618 131546 348854
rect 131782 348618 131866 348854
rect 132102 348618 132134 348854
rect 131514 313174 132134 348618
rect 131514 312938 131546 313174
rect 131782 312938 131866 313174
rect 132102 312938 132134 313174
rect 131514 312854 132134 312938
rect 131514 312618 131546 312854
rect 131782 312618 131866 312854
rect 132102 312618 132134 312854
rect 131514 285308 132134 312618
rect 135234 352894 135854 378000
rect 136035 377980 136036 378044
rect 136100 377980 136101 378044
rect 136035 377979 136101 377980
rect 138611 378044 138677 378045
rect 138611 377980 138612 378044
rect 138676 377980 138677 378044
rect 141003 378044 141069 378045
rect 138611 377979 138677 377980
rect 135234 352658 135266 352894
rect 135502 352658 135586 352894
rect 135822 352658 135854 352894
rect 135234 352574 135854 352658
rect 135234 352338 135266 352574
rect 135502 352338 135586 352574
rect 135822 352338 135854 352574
rect 135234 316894 135854 352338
rect 135234 316658 135266 316894
rect 135502 316658 135586 316894
rect 135822 316658 135854 316894
rect 135234 316574 135854 316658
rect 135234 316338 135266 316574
rect 135502 316338 135586 316574
rect 135822 316338 135854 316574
rect 133459 285700 133525 285701
rect 133459 285636 133460 285700
rect 133524 285636 133525 285700
rect 133459 285635 133525 285636
rect 128675 285156 128741 285157
rect 128675 285092 128676 285156
rect 128740 285092 128741 285156
rect 128675 285091 128741 285092
rect 131067 285156 131133 285157
rect 131067 285092 131068 285156
rect 131132 285092 131133 285156
rect 131067 285091 131133 285092
rect 128678 283930 128738 285091
rect 131070 283930 131130 285091
rect 120766 283870 121060 283930
rect 123526 283870 123644 283930
rect 110936 283220 110996 283870
rect 113656 283220 113716 283870
rect 116104 283220 116164 283870
rect 118552 283220 118612 283870
rect 121000 283220 121060 283870
rect 123584 283220 123644 283870
rect 125896 283870 125978 283930
rect 128616 283870 128738 283930
rect 131064 283870 131130 283930
rect 133462 283930 133522 285635
rect 135234 285308 135854 316338
rect 138954 356614 139574 378000
rect 141003 377980 141004 378044
rect 141068 377980 141069 378044
rect 141003 377979 141069 377980
rect 143395 378044 143461 378045
rect 143395 377980 143396 378044
rect 143460 377980 143461 378044
rect 143395 377979 143461 377980
rect 138954 356378 138986 356614
rect 139222 356378 139306 356614
rect 139542 356378 139574 356614
rect 138954 356294 139574 356378
rect 138954 356058 138986 356294
rect 139222 356058 139306 356294
rect 139542 356058 139574 356294
rect 138954 320614 139574 356058
rect 138954 320378 138986 320614
rect 139222 320378 139306 320614
rect 139542 320378 139574 320614
rect 138954 320294 139574 320378
rect 138954 320058 138986 320294
rect 139222 320058 139306 320294
rect 139542 320058 139574 320294
rect 136035 286244 136101 286245
rect 136035 286180 136036 286244
rect 136100 286180 136101 286244
rect 136035 286179 136101 286180
rect 138427 286244 138493 286245
rect 138427 286180 138428 286244
rect 138492 286180 138493 286244
rect 138427 286179 138493 286180
rect 136038 283930 136098 286179
rect 138430 283930 138490 286179
rect 138954 285308 139574 320058
rect 145794 363454 146414 378000
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 145794 327454 146414 362898
rect 145794 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 146414 327454
rect 145794 327134 146414 327218
rect 145794 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 146414 327134
rect 145794 291454 146414 326898
rect 145794 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 146414 291454
rect 145794 291134 146414 291218
rect 145794 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 146414 291134
rect 143579 286244 143645 286245
rect 143579 286180 143580 286244
rect 143644 286180 143645 286244
rect 143579 286179 143645 286180
rect 141003 285700 141069 285701
rect 141003 285636 141004 285700
rect 141068 285636 141069 285700
rect 141003 285635 141069 285636
rect 141006 283930 141066 285635
rect 143582 283930 143642 286179
rect 145794 285308 146414 290898
rect 149514 367174 150134 378000
rect 149514 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 150134 367174
rect 149514 366854 150134 366938
rect 149514 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 150134 366854
rect 149514 331174 150134 366618
rect 149514 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 150134 331174
rect 149514 330854 150134 330938
rect 149514 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 150134 330854
rect 149514 295174 150134 330618
rect 149514 294938 149546 295174
rect 149782 294938 149866 295174
rect 150102 294938 150134 295174
rect 149514 294854 150134 294938
rect 149514 294618 149546 294854
rect 149782 294618 149866 294854
rect 150102 294618 150134 294854
rect 149514 285308 150134 294618
rect 153234 370894 153854 378000
rect 153234 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 153854 370894
rect 153234 370574 153854 370658
rect 153234 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 153854 370574
rect 153234 334894 153854 370338
rect 153234 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 153854 334894
rect 153234 334574 153854 334658
rect 153234 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 153854 334574
rect 153234 298894 153854 334338
rect 153234 298658 153266 298894
rect 153502 298658 153586 298894
rect 153822 298658 153854 298894
rect 153234 298574 153854 298658
rect 153234 298338 153266 298574
rect 153502 298338 153586 298574
rect 153822 298338 153854 298574
rect 151123 285700 151189 285701
rect 151123 285636 151124 285700
rect 151188 285636 151189 285700
rect 151123 285635 151189 285636
rect 148547 284884 148613 284885
rect 148547 284820 148548 284884
rect 148612 284820 148613 284884
rect 148547 284819 148613 284820
rect 145971 284748 146037 284749
rect 145971 284684 145972 284748
rect 146036 284684 146037 284748
rect 145971 284683 146037 284684
rect 133462 283870 133572 283930
rect 125896 283220 125956 283870
rect 128616 283220 128676 283870
rect 131064 283220 131124 283870
rect 133512 283220 133572 283870
rect 135960 283870 136098 283930
rect 138408 283870 138490 283930
rect 140992 283870 141066 283930
rect 143576 283870 143642 283930
rect 145974 283930 146034 284683
rect 148550 283930 148610 284819
rect 151126 283930 151186 285635
rect 153234 285308 153854 298338
rect 156954 374614 157574 378000
rect 156954 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 157574 374614
rect 156954 374294 157574 374378
rect 156954 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 157574 374294
rect 156954 338614 157574 374058
rect 156954 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 157574 338614
rect 156954 338294 157574 338378
rect 156954 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 157574 338294
rect 156954 302614 157574 338058
rect 156954 302378 156986 302614
rect 157222 302378 157306 302614
rect 157542 302378 157574 302614
rect 156954 302294 157574 302378
rect 156954 302058 156986 302294
rect 157222 302058 157306 302294
rect 157542 302058 157574 302294
rect 154067 285700 154133 285701
rect 154067 285636 154068 285700
rect 154132 285636 154133 285700
rect 154067 285635 154133 285636
rect 156091 285700 156157 285701
rect 156091 285636 156092 285700
rect 156156 285636 156157 285700
rect 156091 285635 156157 285636
rect 154070 283930 154130 285635
rect 156094 283930 156154 285635
rect 156954 285308 157574 302058
rect 163794 345454 164414 378000
rect 163794 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 164414 345454
rect 163794 345134 164414 345218
rect 163794 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 164414 345134
rect 163794 309454 164414 344898
rect 163794 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 164414 309454
rect 163794 309134 164414 309218
rect 163794 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 164414 309134
rect 163794 285308 164414 308898
rect 167514 349174 168134 378000
rect 167514 348938 167546 349174
rect 167782 348938 167866 349174
rect 168102 348938 168134 349174
rect 167514 348854 168134 348938
rect 167514 348618 167546 348854
rect 167782 348618 167866 348854
rect 168102 348618 168134 348854
rect 167514 313174 168134 348618
rect 167514 312938 167546 313174
rect 167782 312938 167866 313174
rect 168102 312938 168134 313174
rect 167514 312854 168134 312938
rect 167514 312618 167546 312854
rect 167782 312618 167866 312854
rect 168102 312618 168134 312854
rect 167514 285308 168134 312618
rect 171234 352894 171854 378000
rect 173206 376957 173266 379750
rect 173390 377093 173450 379750
rect 173387 377092 173453 377093
rect 173387 377028 173388 377092
rect 173452 377028 173453 377092
rect 173387 377027 173453 377028
rect 173203 376956 173269 376957
rect 173203 376892 173204 376956
rect 173268 376892 173269 376956
rect 173203 376891 173269 376892
rect 171234 352658 171266 352894
rect 171502 352658 171586 352894
rect 171822 352658 171854 352894
rect 171234 352574 171854 352658
rect 171234 352338 171266 352574
rect 171502 352338 171586 352574
rect 171822 352338 171854 352574
rect 171234 316894 171854 352338
rect 171234 316658 171266 316894
rect 171502 316658 171586 316894
rect 171822 316658 171854 316894
rect 171234 316574 171854 316658
rect 171234 316338 171266 316574
rect 171502 316338 171586 316574
rect 171822 316338 171854 316574
rect 169707 286244 169773 286245
rect 169707 286180 169708 286244
rect 169772 286180 169773 286244
rect 169707 286179 169773 286180
rect 168419 285700 168485 285701
rect 168419 285636 168420 285700
rect 168484 285636 168485 285700
rect 168419 285635 168485 285636
rect 145974 283870 146084 283930
rect 135960 283220 136020 283870
rect 138408 283220 138468 283870
rect 140992 283220 141052 283870
rect 143576 283220 143636 283870
rect 146024 283220 146084 283870
rect 148472 283870 148610 283930
rect 151056 283870 151186 283930
rect 153368 283870 154130 283930
rect 156088 283870 156154 283930
rect 168422 283930 168482 285635
rect 169710 283930 169770 286179
rect 171234 285308 171854 316338
rect 174954 356614 175574 378000
rect 174954 356378 174986 356614
rect 175222 356378 175306 356614
rect 175542 356378 175574 356614
rect 174954 356294 175574 356378
rect 174954 356058 174986 356294
rect 175222 356058 175306 356294
rect 175542 356058 175574 356294
rect 174954 320614 175574 356058
rect 174954 320378 174986 320614
rect 175222 320378 175306 320614
rect 175542 320378 175574 320614
rect 174954 320294 175574 320378
rect 174954 320058 174986 320294
rect 175222 320058 175306 320294
rect 175542 320058 175574 320294
rect 174954 285308 175574 320058
rect 181794 363454 182414 378000
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 181794 327454 182414 362898
rect 181794 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 182414 327454
rect 181794 327134 182414 327218
rect 181794 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 182414 327134
rect 181794 291454 182414 326898
rect 181794 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 182414 291454
rect 181794 291134 182414 291218
rect 181794 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 182414 291134
rect 181794 285308 182414 290898
rect 185514 367174 186134 378000
rect 185514 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 186134 367174
rect 185514 366854 186134 366938
rect 185514 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 186134 366854
rect 185514 331174 186134 366618
rect 185514 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 186134 331174
rect 185514 330854 186134 330938
rect 185514 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 186134 330854
rect 185514 295174 186134 330618
rect 185514 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 186134 295174
rect 185514 294854 186134 294938
rect 185514 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 186134 294854
rect 185514 285308 186134 294618
rect 189234 370894 189854 406338
rect 189234 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 189854 370894
rect 189234 370574 189854 370658
rect 189234 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 189854 370574
rect 189234 334894 189854 370338
rect 189234 334658 189266 334894
rect 189502 334658 189586 334894
rect 189822 334658 189854 334894
rect 189234 334574 189854 334658
rect 189234 334338 189266 334574
rect 189502 334338 189586 334574
rect 189822 334338 189854 334574
rect 189234 298894 189854 334338
rect 189234 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 189854 298894
rect 189234 298574 189854 298658
rect 189234 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 189854 298574
rect 187187 285972 187253 285973
rect 187187 285908 187188 285972
rect 187252 285908 187253 285972
rect 187187 285907 187253 285908
rect 180747 284068 180813 284069
rect 180747 284004 180748 284068
rect 180812 284004 180813 284068
rect 180747 284003 180813 284004
rect 168422 283870 168524 283930
rect 148472 283220 148532 283870
rect 151056 283220 151116 283870
rect 153368 283220 153428 283870
rect 156088 283220 156148 283870
rect 168464 283220 168524 283870
rect 169688 283870 169770 283930
rect 180750 283930 180810 284003
rect 180750 283870 180900 283930
rect 169688 283220 169748 283870
rect 180840 283220 180900 283870
rect 186819 277540 186885 277541
rect 186819 277476 186820 277540
rect 186884 277476 186885 277540
rect 186819 277475 186885 277476
rect 50272 273454 50620 273486
rect 50272 273218 50328 273454
rect 50564 273218 50620 273454
rect 50272 273134 50620 273218
rect 50272 272898 50328 273134
rect 50564 272898 50620 273134
rect 50272 272866 50620 272898
rect 186000 273454 186348 273486
rect 186000 273218 186056 273454
rect 186292 273218 186348 273454
rect 186000 273134 186348 273218
rect 186000 272898 186056 273134
rect 186292 272898 186348 273134
rect 186000 272866 186348 272898
rect 45234 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 45854 262894
rect 45234 262574 45854 262658
rect 45234 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 45854 262574
rect 45234 226894 45854 262338
rect 50952 255454 51300 255486
rect 50952 255218 51008 255454
rect 51244 255218 51300 255454
rect 50952 255134 51300 255218
rect 50952 254898 51008 255134
rect 51244 254898 51300 255134
rect 50952 254866 51300 254898
rect 185320 255454 185668 255486
rect 185320 255218 185376 255454
rect 185612 255218 185668 255454
rect 185320 255134 185668 255218
rect 185320 254898 185376 255134
rect 185612 254898 185668 255134
rect 185320 254866 185668 254898
rect 50272 237454 50620 237486
rect 50272 237218 50328 237454
rect 50564 237218 50620 237454
rect 50272 237134 50620 237218
rect 50272 236898 50328 237134
rect 50564 236898 50620 237134
rect 50272 236866 50620 236898
rect 186000 237454 186348 237486
rect 186000 237218 186056 237454
rect 186292 237218 186348 237454
rect 186000 237134 186348 237218
rect 186000 236898 186056 237134
rect 186292 236898 186348 237134
rect 186000 236866 186348 236898
rect 45234 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 45854 226894
rect 45234 226574 45854 226658
rect 45234 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 45854 226574
rect 45234 190894 45854 226338
rect 50952 219454 51300 219486
rect 50952 219218 51008 219454
rect 51244 219218 51300 219454
rect 50952 219134 51300 219218
rect 50952 218898 51008 219134
rect 51244 218898 51300 219134
rect 50952 218866 51300 218898
rect 185320 219454 185668 219486
rect 185320 219218 185376 219454
rect 185612 219218 185668 219454
rect 185320 219134 185668 219218
rect 185320 218898 185376 219134
rect 185612 218898 185668 219134
rect 185320 218866 185668 218898
rect 50272 201454 50620 201486
rect 50272 201218 50328 201454
rect 50564 201218 50620 201454
rect 50272 201134 50620 201218
rect 50272 200898 50328 201134
rect 50564 200898 50620 201134
rect 50272 200866 50620 200898
rect 186000 201454 186348 201486
rect 186000 201218 186056 201454
rect 186292 201218 186348 201454
rect 186000 201134 186348 201218
rect 186000 200898 186056 201134
rect 186292 200898 186348 201134
rect 186000 200866 186348 200898
rect 66056 199610 66116 200130
rect 67144 199610 67204 200130
rect 68232 199610 68292 200130
rect 69592 199610 69652 200130
rect 70544 199610 70604 200130
rect 66056 199550 66178 199610
rect 67144 199550 67282 199610
rect 68232 199550 68386 199610
rect 69592 199550 69674 199610
rect 45234 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 45854 190894
rect 45234 190574 45854 190658
rect 45234 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 45854 190574
rect 45234 154894 45854 190338
rect 45234 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 45854 154894
rect 45234 154574 45854 154658
rect 45234 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 45854 154574
rect 45234 118894 45854 154338
rect 45234 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 45854 118894
rect 45234 118574 45854 118658
rect 45234 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 45854 118574
rect 45234 82894 45854 118338
rect 45234 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 45854 82894
rect 45234 82574 45854 82658
rect 45234 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 45854 82574
rect 45234 46894 45854 82338
rect 45234 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 45854 46894
rect 45234 46574 45854 46658
rect 45234 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 45854 46574
rect 45234 10894 45854 46338
rect 45234 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 45854 10894
rect 45234 10574 45854 10658
rect 45234 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 45854 10574
rect 45234 -4186 45854 10338
rect 45234 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 45854 -4186
rect 45234 -4506 45854 -4422
rect 45234 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 45854 -4506
rect 45234 -5734 45854 -4742
rect 48954 194614 49574 198000
rect 48954 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 49574 194614
rect 48954 194294 49574 194378
rect 48954 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 49574 194294
rect 48954 158614 49574 194058
rect 48954 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 49574 158614
rect 48954 158294 49574 158378
rect 48954 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 49574 158294
rect 48954 122614 49574 158058
rect 48954 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 49574 122614
rect 48954 122294 49574 122378
rect 48954 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 49574 122294
rect 48954 86614 49574 122058
rect 48954 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 49574 86614
rect 48954 86294 49574 86378
rect 48954 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 49574 86294
rect 48954 50614 49574 86058
rect 48954 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 49574 50614
rect 48954 50294 49574 50378
rect 48954 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 49574 50294
rect 48954 14614 49574 50058
rect 48954 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 49574 14614
rect 48954 14294 49574 14378
rect 48954 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 49574 14294
rect 30954 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 31574 -7066
rect 30954 -7386 31574 -7302
rect 30954 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 31574 -7386
rect 30954 -7654 31574 -7622
rect 48954 -6106 49574 14058
rect 55794 165454 56414 198000
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -1306 56414 20898
rect 55794 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 56414 -1306
rect 55794 -1626 56414 -1542
rect 55794 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 56414 -1626
rect 55794 -1894 56414 -1862
rect 59514 169174 60134 198000
rect 59514 168938 59546 169174
rect 59782 168938 59866 169174
rect 60102 168938 60134 169174
rect 59514 168854 60134 168938
rect 59514 168618 59546 168854
rect 59782 168618 59866 168854
rect 60102 168618 60134 168854
rect 59514 133174 60134 168618
rect 59514 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 60134 133174
rect 59514 132854 60134 132938
rect 59514 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 60134 132854
rect 59514 97174 60134 132618
rect 59514 96938 59546 97174
rect 59782 96938 59866 97174
rect 60102 96938 60134 97174
rect 59514 96854 60134 96938
rect 59514 96618 59546 96854
rect 59782 96618 59866 96854
rect 60102 96618 60134 96854
rect 59514 61174 60134 96618
rect 59514 60938 59546 61174
rect 59782 60938 59866 61174
rect 60102 60938 60134 61174
rect 59514 60854 60134 60938
rect 59514 60618 59546 60854
rect 59782 60618 59866 60854
rect 60102 60618 60134 60854
rect 59514 25174 60134 60618
rect 59514 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 60134 25174
rect 59514 24854 60134 24938
rect 59514 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 60134 24854
rect 59514 -3226 60134 24618
rect 59514 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 60134 -3226
rect 59514 -3546 60134 -3462
rect 59514 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 60134 -3546
rect 59514 -3814 60134 -3782
rect 63234 172894 63854 198000
rect 66118 197437 66178 199550
rect 67222 198253 67282 199550
rect 67219 198252 67285 198253
rect 67219 198188 67220 198252
rect 67284 198188 67285 198252
rect 67219 198187 67285 198188
rect 66115 197436 66181 197437
rect 66115 197372 66116 197436
rect 66180 197372 66181 197436
rect 66115 197371 66181 197372
rect 63234 172658 63266 172894
rect 63502 172658 63586 172894
rect 63822 172658 63854 172894
rect 63234 172574 63854 172658
rect 63234 172338 63266 172574
rect 63502 172338 63586 172574
rect 63822 172338 63854 172574
rect 63234 136894 63854 172338
rect 63234 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 63854 136894
rect 63234 136574 63854 136658
rect 63234 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 63854 136574
rect 63234 100894 63854 136338
rect 63234 100658 63266 100894
rect 63502 100658 63586 100894
rect 63822 100658 63854 100894
rect 63234 100574 63854 100658
rect 63234 100338 63266 100574
rect 63502 100338 63586 100574
rect 63822 100338 63854 100574
rect 63234 64894 63854 100338
rect 63234 64658 63266 64894
rect 63502 64658 63586 64894
rect 63822 64658 63854 64894
rect 63234 64574 63854 64658
rect 63234 64338 63266 64574
rect 63502 64338 63586 64574
rect 63822 64338 63854 64574
rect 63234 28894 63854 64338
rect 63234 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 63854 28894
rect 63234 28574 63854 28658
rect 63234 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 63854 28574
rect 63234 -5146 63854 28338
rect 63234 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 63854 -5146
rect 63234 -5466 63854 -5382
rect 63234 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 63854 -5466
rect 63234 -5734 63854 -5702
rect 66954 176614 67574 198000
rect 68326 197437 68386 199550
rect 69614 197437 69674 199550
rect 70534 199550 70604 199610
rect 71768 199610 71828 200130
rect 73128 199610 73188 200130
rect 71768 199550 71882 199610
rect 70534 198661 70594 199550
rect 71822 199477 71882 199550
rect 73110 199550 73188 199610
rect 74214 200070 74276 200130
rect 71819 199476 71885 199477
rect 71819 199412 71820 199476
rect 71884 199412 71885 199476
rect 71819 199411 71885 199412
rect 70531 198660 70597 198661
rect 70531 198596 70532 198660
rect 70596 198596 70597 198660
rect 70531 198595 70597 198596
rect 73110 197437 73170 199550
rect 74214 198253 74274 200070
rect 75440 199610 75500 200130
rect 76528 199610 76588 200130
rect 77616 199610 77676 200130
rect 78296 199610 78356 200130
rect 75440 199550 75562 199610
rect 76528 199550 76666 199610
rect 77616 199550 77770 199610
rect 74211 198252 74277 198253
rect 74211 198188 74212 198252
rect 74276 198188 74277 198252
rect 74211 198187 74277 198188
rect 75502 198117 75562 199550
rect 76606 198661 76666 199550
rect 77710 199477 77770 199550
rect 78262 199550 78356 199610
rect 78704 199610 78764 200130
rect 80064 199610 80124 200130
rect 80744 199610 80804 200130
rect 81288 199610 81348 200130
rect 82376 199610 82436 200130
rect 83464 199610 83524 200130
rect 78704 199550 78874 199610
rect 80064 199550 80162 199610
rect 80744 199550 80898 199610
rect 81288 199550 81450 199610
rect 82376 199550 82554 199610
rect 77707 199476 77773 199477
rect 77707 199412 77708 199476
rect 77772 199412 77773 199476
rect 77707 199411 77773 199412
rect 76603 198660 76669 198661
rect 76603 198596 76604 198660
rect 76668 198596 76669 198660
rect 76603 198595 76669 198596
rect 75499 198116 75565 198117
rect 75499 198052 75500 198116
rect 75564 198052 75565 198116
rect 75499 198051 75565 198052
rect 68323 197436 68389 197437
rect 68323 197372 68324 197436
rect 68388 197372 68389 197436
rect 68323 197371 68389 197372
rect 69611 197436 69677 197437
rect 69611 197372 69612 197436
rect 69676 197372 69677 197436
rect 69611 197371 69677 197372
rect 73107 197436 73173 197437
rect 73107 197372 73108 197436
rect 73172 197372 73173 197436
rect 73107 197371 73173 197372
rect 66954 176378 66986 176614
rect 67222 176378 67306 176614
rect 67542 176378 67574 176614
rect 66954 176294 67574 176378
rect 66954 176058 66986 176294
rect 67222 176058 67306 176294
rect 67542 176058 67574 176294
rect 66954 140614 67574 176058
rect 66954 140378 66986 140614
rect 67222 140378 67306 140614
rect 67542 140378 67574 140614
rect 66954 140294 67574 140378
rect 66954 140058 66986 140294
rect 67222 140058 67306 140294
rect 67542 140058 67574 140294
rect 66954 104614 67574 140058
rect 66954 104378 66986 104614
rect 67222 104378 67306 104614
rect 67542 104378 67574 104614
rect 66954 104294 67574 104378
rect 66954 104058 66986 104294
rect 67222 104058 67306 104294
rect 67542 104058 67574 104294
rect 66954 68614 67574 104058
rect 66954 68378 66986 68614
rect 67222 68378 67306 68614
rect 67542 68378 67574 68614
rect 66954 68294 67574 68378
rect 66954 68058 66986 68294
rect 67222 68058 67306 68294
rect 67542 68058 67574 68294
rect 66954 32614 67574 68058
rect 66954 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 67574 32614
rect 66954 32294 67574 32378
rect 66954 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 67574 32294
rect 48954 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 49574 -6106
rect 48954 -6426 49574 -6342
rect 48954 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 49574 -6426
rect 48954 -7654 49574 -6662
rect 66954 -7066 67574 32058
rect 73794 183454 74414 198000
rect 73794 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 74414 183454
rect 73794 183134 74414 183218
rect 73794 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 74414 183134
rect 73794 147454 74414 182898
rect 73794 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 74414 147454
rect 73794 147134 74414 147218
rect 73794 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 74414 147134
rect 73794 111454 74414 146898
rect 73794 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 74414 111454
rect 73794 111134 74414 111218
rect 73794 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 74414 111134
rect 73794 75454 74414 110898
rect 73794 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 74414 75454
rect 73794 75134 74414 75218
rect 73794 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 74414 75134
rect 73794 39454 74414 74898
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -1894 74414 -902
rect 77514 187174 78134 198000
rect 78262 197437 78322 199550
rect 78814 198661 78874 199550
rect 80102 198661 80162 199550
rect 78811 198660 78877 198661
rect 78811 198596 78812 198660
rect 78876 198596 78877 198660
rect 78811 198595 78877 198596
rect 80099 198660 80165 198661
rect 80099 198596 80100 198660
rect 80164 198596 80165 198660
rect 80099 198595 80165 198596
rect 80838 197437 80898 199550
rect 81390 199477 81450 199550
rect 82494 199477 82554 199550
rect 83414 199550 83524 199610
rect 83598 200070 83660 200130
rect 83414 199477 83474 199550
rect 81387 199476 81453 199477
rect 81387 199412 81388 199476
rect 81452 199412 81453 199476
rect 81387 199411 81453 199412
rect 82491 199476 82557 199477
rect 82491 199412 82492 199476
rect 82556 199412 82557 199476
rect 82491 199411 82557 199412
rect 83411 199476 83477 199477
rect 83411 199412 83412 199476
rect 83476 199412 83477 199476
rect 83411 199411 83477 199412
rect 78259 197436 78325 197437
rect 78259 197372 78260 197436
rect 78324 197372 78325 197436
rect 78259 197371 78325 197372
rect 80835 197436 80901 197437
rect 80835 197372 80836 197436
rect 80900 197372 80901 197436
rect 80835 197371 80901 197372
rect 77514 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 78134 187174
rect 77514 186854 78134 186938
rect 77514 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 78134 186854
rect 77514 151174 78134 186618
rect 77514 150938 77546 151174
rect 77782 150938 77866 151174
rect 78102 150938 78134 151174
rect 77514 150854 78134 150938
rect 77514 150618 77546 150854
rect 77782 150618 77866 150854
rect 78102 150618 78134 150854
rect 77514 115174 78134 150618
rect 77514 114938 77546 115174
rect 77782 114938 77866 115174
rect 78102 114938 78134 115174
rect 77514 114854 78134 114938
rect 77514 114618 77546 114854
rect 77782 114618 77866 114854
rect 78102 114618 78134 114854
rect 77514 79174 78134 114618
rect 77514 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 78134 79174
rect 77514 78854 78134 78938
rect 77514 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 78134 78854
rect 77514 43174 78134 78618
rect 77514 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 78134 43174
rect 77514 42854 78134 42938
rect 77514 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 78134 42854
rect 77514 7174 78134 42618
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -2266 78134 6618
rect 77514 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 78134 -2266
rect 77514 -2586 78134 -2502
rect 77514 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 78134 -2586
rect 77514 -3814 78134 -2822
rect 81234 190894 81854 198000
rect 83598 197981 83658 200070
rect 84552 199610 84612 200130
rect 85912 199610 85972 200130
rect 84518 199550 84612 199610
rect 85806 199550 85972 199610
rect 86048 199610 86108 200130
rect 87000 199610 87060 200130
rect 88088 199610 88148 200130
rect 88496 199610 88556 200130
rect 89448 199610 89508 200130
rect 90672 199610 90732 200130
rect 91080 199610 91140 200130
rect 91760 199610 91820 200130
rect 92848 199610 92908 200130
rect 93528 200070 93594 200130
rect 86048 199550 86234 199610
rect 87000 199550 87154 199610
rect 88088 199550 88258 199610
rect 88496 199550 88626 199610
rect 89448 199550 89546 199610
rect 90672 199550 90834 199610
rect 91080 199550 91202 199610
rect 91760 199550 91938 199610
rect 84518 198661 84578 199550
rect 84515 198660 84581 198661
rect 84515 198596 84516 198660
rect 84580 198596 84581 198660
rect 84515 198595 84581 198596
rect 85806 198525 85866 199550
rect 86174 199477 86234 199550
rect 86171 199476 86237 199477
rect 86171 199412 86172 199476
rect 86236 199412 86237 199476
rect 86171 199411 86237 199412
rect 87094 198525 87154 199550
rect 88198 198661 88258 199550
rect 88566 198661 88626 199550
rect 88195 198660 88261 198661
rect 88195 198596 88196 198660
rect 88260 198596 88261 198660
rect 88195 198595 88261 198596
rect 88563 198660 88629 198661
rect 88563 198596 88564 198660
rect 88628 198596 88629 198660
rect 88563 198595 88629 198596
rect 85803 198524 85869 198525
rect 85803 198460 85804 198524
rect 85868 198460 85869 198524
rect 85803 198459 85869 198460
rect 87091 198524 87157 198525
rect 87091 198460 87092 198524
rect 87156 198460 87157 198524
rect 87091 198459 87157 198460
rect 89486 198389 89546 199550
rect 90774 198525 90834 199550
rect 91142 198661 91202 199550
rect 91139 198660 91205 198661
rect 91139 198596 91140 198660
rect 91204 198596 91205 198660
rect 91139 198595 91205 198596
rect 90771 198524 90837 198525
rect 90771 198460 90772 198524
rect 90836 198460 90837 198524
rect 90771 198459 90837 198460
rect 89483 198388 89549 198389
rect 89483 198324 89484 198388
rect 89548 198324 89549 198388
rect 89483 198323 89549 198324
rect 91878 198253 91938 199550
rect 92798 199550 92908 199610
rect 92798 198389 92858 199550
rect 93534 198661 93594 200070
rect 93936 199610 93996 200130
rect 93902 199550 93996 199610
rect 95296 199610 95356 200130
rect 95976 199610 96036 200130
rect 95296 199550 95434 199610
rect 93902 198661 93962 199550
rect 93531 198660 93597 198661
rect 93531 198596 93532 198660
rect 93596 198596 93597 198660
rect 93531 198595 93597 198596
rect 93899 198660 93965 198661
rect 93899 198596 93900 198660
rect 93964 198596 93965 198660
rect 93899 198595 93965 198596
rect 95374 198389 95434 199550
rect 95926 199550 96036 199610
rect 96384 199610 96444 200130
rect 97608 199610 97668 200130
rect 96384 199550 96538 199610
rect 95926 198661 95986 199550
rect 95923 198660 95989 198661
rect 95923 198596 95924 198660
rect 95988 198596 95989 198660
rect 95923 198595 95989 198596
rect 96478 198525 96538 199550
rect 97582 199550 97668 199610
rect 98288 199610 98348 200130
rect 98696 199610 98756 200130
rect 99784 200070 99850 200130
rect 98288 199550 98378 199610
rect 96475 198524 96541 198525
rect 96475 198460 96476 198524
rect 96540 198460 96541 198524
rect 96475 198459 96541 198460
rect 92795 198388 92861 198389
rect 92795 198324 92796 198388
rect 92860 198324 92861 198388
rect 92795 198323 92861 198324
rect 95371 198388 95437 198389
rect 95371 198324 95372 198388
rect 95436 198324 95437 198388
rect 95371 198323 95437 198324
rect 91875 198252 91941 198253
rect 91875 198188 91876 198252
rect 91940 198188 91941 198252
rect 91875 198187 91941 198188
rect 83595 197980 83661 197981
rect 83595 197916 83596 197980
rect 83660 197916 83661 197980
rect 83595 197915 83661 197916
rect 81234 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 81854 190894
rect 81234 190574 81854 190658
rect 81234 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 81854 190574
rect 81234 154894 81854 190338
rect 81234 154658 81266 154894
rect 81502 154658 81586 154894
rect 81822 154658 81854 154894
rect 81234 154574 81854 154658
rect 81234 154338 81266 154574
rect 81502 154338 81586 154574
rect 81822 154338 81854 154574
rect 81234 118894 81854 154338
rect 81234 118658 81266 118894
rect 81502 118658 81586 118894
rect 81822 118658 81854 118894
rect 81234 118574 81854 118658
rect 81234 118338 81266 118574
rect 81502 118338 81586 118574
rect 81822 118338 81854 118574
rect 81234 82894 81854 118338
rect 81234 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 81854 82894
rect 81234 82574 81854 82658
rect 81234 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 81854 82574
rect 81234 46894 81854 82338
rect 81234 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 81854 46894
rect 81234 46574 81854 46658
rect 81234 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 81854 46574
rect 81234 10894 81854 46338
rect 81234 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 81854 10894
rect 81234 10574 81854 10658
rect 81234 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 81854 10574
rect 81234 -4186 81854 10338
rect 81234 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 81854 -4186
rect 81234 -4506 81854 -4422
rect 81234 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 81854 -4506
rect 81234 -5734 81854 -4742
rect 84954 194614 85574 198000
rect 84954 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 85574 194614
rect 84954 194294 85574 194378
rect 84954 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 85574 194294
rect 84954 158614 85574 194058
rect 84954 158378 84986 158614
rect 85222 158378 85306 158614
rect 85542 158378 85574 158614
rect 84954 158294 85574 158378
rect 84954 158058 84986 158294
rect 85222 158058 85306 158294
rect 85542 158058 85574 158294
rect 84954 122614 85574 158058
rect 84954 122378 84986 122614
rect 85222 122378 85306 122614
rect 85542 122378 85574 122614
rect 84954 122294 85574 122378
rect 84954 122058 84986 122294
rect 85222 122058 85306 122294
rect 85542 122058 85574 122294
rect 84954 86614 85574 122058
rect 84954 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 85574 86614
rect 84954 86294 85574 86378
rect 84954 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 85574 86294
rect 84954 50614 85574 86058
rect 84954 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 85574 50614
rect 84954 50294 85574 50378
rect 84954 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 85574 50294
rect 84954 14614 85574 50058
rect 84954 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 85574 14614
rect 84954 14294 85574 14378
rect 84954 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 85574 14294
rect 66954 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 67574 -7066
rect 66954 -7386 67574 -7302
rect 66954 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 67574 -7386
rect 66954 -7654 67574 -7622
rect 84954 -6106 85574 14058
rect 91794 165454 92414 198000
rect 91794 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 92414 165454
rect 91794 165134 92414 165218
rect 91794 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 92414 165134
rect 91794 129454 92414 164898
rect 91794 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 92414 129454
rect 91794 129134 92414 129218
rect 91794 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 92414 129134
rect 91794 93454 92414 128898
rect 91794 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 92414 93454
rect 91794 93134 92414 93218
rect 91794 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 92414 93134
rect 91794 57454 92414 92898
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -1306 92414 20898
rect 91794 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 92414 -1306
rect 91794 -1626 92414 -1542
rect 91794 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 92414 -1626
rect 91794 -1894 92414 -1862
rect 95514 169174 96134 198000
rect 97582 197437 97642 199550
rect 98318 198661 98378 199550
rect 98686 199550 98756 199610
rect 98315 198660 98381 198661
rect 98315 198596 98316 198660
rect 98380 198596 98381 198660
rect 98315 198595 98381 198596
rect 98686 197573 98746 199550
rect 99790 198661 99850 200070
rect 101008 199610 101068 200130
rect 100894 199550 101068 199610
rect 101144 199610 101204 200130
rect 102232 199610 102292 200130
rect 103320 199610 103380 200130
rect 101144 199550 101322 199610
rect 100894 198661 100954 199550
rect 99787 198660 99853 198661
rect 99787 198596 99788 198660
rect 99852 198596 99853 198660
rect 99787 198595 99853 198596
rect 100891 198660 100957 198661
rect 100891 198596 100892 198660
rect 100956 198596 100957 198660
rect 100891 198595 100957 198596
rect 101262 198253 101322 199550
rect 102182 199550 102292 199610
rect 103286 199550 103380 199610
rect 103592 199610 103652 200130
rect 104408 199610 104468 200130
rect 103592 199550 103714 199610
rect 102182 198661 102242 199550
rect 103286 198933 103346 199550
rect 103654 199477 103714 199550
rect 104390 199550 104468 199610
rect 105768 199610 105828 200130
rect 106040 200070 106106 200130
rect 105768 199550 105922 199610
rect 103651 199476 103717 199477
rect 103651 199412 103652 199476
rect 103716 199412 103717 199476
rect 103651 199411 103717 199412
rect 103283 198932 103349 198933
rect 103283 198868 103284 198932
rect 103348 198868 103349 198932
rect 103283 198867 103349 198868
rect 102179 198660 102245 198661
rect 102179 198596 102180 198660
rect 102244 198596 102245 198660
rect 102179 198595 102245 198596
rect 101259 198252 101325 198253
rect 101259 198188 101260 198252
rect 101324 198188 101325 198252
rect 101259 198187 101325 198188
rect 104390 198117 104450 199550
rect 104387 198116 104453 198117
rect 104387 198052 104388 198116
rect 104452 198052 104453 198116
rect 104387 198051 104453 198052
rect 98683 197572 98749 197573
rect 98683 197508 98684 197572
rect 98748 197508 98749 197572
rect 98683 197507 98749 197508
rect 97579 197436 97645 197437
rect 97579 197372 97580 197436
rect 97644 197372 97645 197436
rect 97579 197371 97645 197372
rect 95514 168938 95546 169174
rect 95782 168938 95866 169174
rect 96102 168938 96134 169174
rect 95514 168854 96134 168938
rect 95514 168618 95546 168854
rect 95782 168618 95866 168854
rect 96102 168618 96134 168854
rect 95514 133174 96134 168618
rect 95514 132938 95546 133174
rect 95782 132938 95866 133174
rect 96102 132938 96134 133174
rect 95514 132854 96134 132938
rect 95514 132618 95546 132854
rect 95782 132618 95866 132854
rect 96102 132618 96134 132854
rect 95514 97174 96134 132618
rect 95514 96938 95546 97174
rect 95782 96938 95866 97174
rect 96102 96938 96134 97174
rect 95514 96854 96134 96938
rect 95514 96618 95546 96854
rect 95782 96618 95866 96854
rect 96102 96618 96134 96854
rect 95514 61174 96134 96618
rect 95514 60938 95546 61174
rect 95782 60938 95866 61174
rect 96102 60938 96134 61174
rect 95514 60854 96134 60938
rect 95514 60618 95546 60854
rect 95782 60618 95866 60854
rect 96102 60618 96134 60854
rect 95514 25174 96134 60618
rect 95514 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 96134 25174
rect 95514 24854 96134 24938
rect 95514 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 96134 24854
rect 95514 -3226 96134 24618
rect 95514 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 96134 -3226
rect 95514 -3546 96134 -3462
rect 95514 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 96134 -3546
rect 95514 -3814 96134 -3782
rect 99234 172894 99854 198000
rect 99234 172658 99266 172894
rect 99502 172658 99586 172894
rect 99822 172658 99854 172894
rect 99234 172574 99854 172658
rect 99234 172338 99266 172574
rect 99502 172338 99586 172574
rect 99822 172338 99854 172574
rect 99234 136894 99854 172338
rect 99234 136658 99266 136894
rect 99502 136658 99586 136894
rect 99822 136658 99854 136894
rect 99234 136574 99854 136658
rect 99234 136338 99266 136574
rect 99502 136338 99586 136574
rect 99822 136338 99854 136574
rect 99234 100894 99854 136338
rect 99234 100658 99266 100894
rect 99502 100658 99586 100894
rect 99822 100658 99854 100894
rect 99234 100574 99854 100658
rect 99234 100338 99266 100574
rect 99502 100338 99586 100574
rect 99822 100338 99854 100574
rect 99234 64894 99854 100338
rect 99234 64658 99266 64894
rect 99502 64658 99586 64894
rect 99822 64658 99854 64894
rect 99234 64574 99854 64658
rect 99234 64338 99266 64574
rect 99502 64338 99586 64574
rect 99822 64338 99854 64574
rect 99234 28894 99854 64338
rect 99234 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 99854 28894
rect 99234 28574 99854 28658
rect 99234 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 99854 28574
rect 99234 -5146 99854 28338
rect 99234 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 99854 -5146
rect 99234 -5466 99854 -5382
rect 99234 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 99854 -5466
rect 99234 -5734 99854 -5702
rect 102954 176614 103574 198000
rect 105862 197981 105922 199550
rect 106046 198661 106106 200070
rect 106992 199610 107052 200130
rect 108080 199610 108140 200130
rect 108488 199610 108548 200130
rect 109168 200070 109234 200130
rect 106966 199550 107052 199610
rect 108070 199550 108140 199610
rect 108438 199550 108548 199610
rect 106966 198661 107026 199550
rect 106043 198660 106109 198661
rect 106043 198596 106044 198660
rect 106108 198596 106109 198660
rect 106043 198595 106109 198596
rect 106963 198660 107029 198661
rect 106963 198596 106964 198660
rect 107028 198596 107029 198660
rect 106963 198595 107029 198596
rect 105859 197980 105925 197981
rect 105859 197916 105860 197980
rect 105924 197916 105925 197980
rect 105859 197915 105925 197916
rect 108070 197165 108130 199550
rect 108438 198661 108498 199550
rect 108435 198660 108501 198661
rect 108435 198596 108436 198660
rect 108500 198596 108501 198660
rect 108435 198595 108501 198596
rect 108067 197164 108133 197165
rect 108067 197100 108068 197164
rect 108132 197100 108133 197164
rect 108067 197099 108133 197100
rect 109174 197029 109234 200070
rect 110936 199610 110996 200130
rect 113520 199610 113580 200130
rect 115968 199610 116028 200130
rect 118280 199610 118340 200130
rect 121000 199610 121060 200130
rect 110936 199550 111074 199610
rect 113520 199550 113650 199610
rect 115968 199550 116042 199610
rect 118280 199550 118434 199610
rect 109171 197028 109237 197029
rect 109171 196964 109172 197028
rect 109236 196964 109237 197028
rect 109171 196963 109237 196964
rect 102954 176378 102986 176614
rect 103222 176378 103306 176614
rect 103542 176378 103574 176614
rect 102954 176294 103574 176378
rect 102954 176058 102986 176294
rect 103222 176058 103306 176294
rect 103542 176058 103574 176294
rect 102954 140614 103574 176058
rect 102954 140378 102986 140614
rect 103222 140378 103306 140614
rect 103542 140378 103574 140614
rect 102954 140294 103574 140378
rect 102954 140058 102986 140294
rect 103222 140058 103306 140294
rect 103542 140058 103574 140294
rect 102954 104614 103574 140058
rect 102954 104378 102986 104614
rect 103222 104378 103306 104614
rect 103542 104378 103574 104614
rect 102954 104294 103574 104378
rect 102954 104058 102986 104294
rect 103222 104058 103306 104294
rect 103542 104058 103574 104294
rect 102954 68614 103574 104058
rect 102954 68378 102986 68614
rect 103222 68378 103306 68614
rect 103542 68378 103574 68614
rect 102954 68294 103574 68378
rect 102954 68058 102986 68294
rect 103222 68058 103306 68294
rect 103542 68058 103574 68294
rect 102954 32614 103574 68058
rect 102954 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 103574 32614
rect 102954 32294 103574 32378
rect 102954 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 103574 32294
rect 84954 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 85574 -6106
rect 84954 -6426 85574 -6342
rect 84954 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 85574 -6426
rect 84954 -7654 85574 -6662
rect 102954 -7066 103574 32058
rect 109794 183454 110414 198000
rect 111014 197981 111074 199550
rect 113590 198661 113650 199550
rect 113587 198660 113653 198661
rect 113587 198596 113588 198660
rect 113652 198596 113653 198660
rect 113587 198595 113653 198596
rect 111011 197980 111077 197981
rect 111011 197916 111012 197980
rect 111076 197916 111077 197980
rect 111011 197915 111077 197916
rect 109794 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 110414 183454
rect 109794 183134 110414 183218
rect 109794 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 110414 183134
rect 109794 147454 110414 182898
rect 109794 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 110414 147454
rect 109794 147134 110414 147218
rect 109794 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 110414 147134
rect 109794 111454 110414 146898
rect 109794 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 110414 111454
rect 109794 111134 110414 111218
rect 109794 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 110414 111134
rect 109794 75454 110414 110898
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 109794 39454 110414 74898
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -1894 110414 -902
rect 113514 187174 114134 198000
rect 115982 197845 116042 199550
rect 115979 197844 116045 197845
rect 115979 197780 115980 197844
rect 116044 197780 116045 197844
rect 115979 197779 116045 197780
rect 113514 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 114134 187174
rect 113514 186854 114134 186938
rect 113514 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 114134 186854
rect 113514 151174 114134 186618
rect 113514 150938 113546 151174
rect 113782 150938 113866 151174
rect 114102 150938 114134 151174
rect 113514 150854 114134 150938
rect 113514 150618 113546 150854
rect 113782 150618 113866 150854
rect 114102 150618 114134 150854
rect 113514 115174 114134 150618
rect 113514 114938 113546 115174
rect 113782 114938 113866 115174
rect 114102 114938 114134 115174
rect 113514 114854 114134 114938
rect 113514 114618 113546 114854
rect 113782 114618 113866 114854
rect 114102 114618 114134 114854
rect 113514 79174 114134 114618
rect 113514 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 114134 79174
rect 113514 78854 114134 78938
rect 113514 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 114134 78854
rect 113514 43174 114134 78618
rect 113514 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 114134 43174
rect 113514 42854 114134 42938
rect 113514 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 114134 42854
rect 113514 7174 114134 42618
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 113514 -2266 114134 6618
rect 113514 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 114134 -2266
rect 113514 -2586 114134 -2502
rect 113514 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 114134 -2586
rect 113514 -3814 114134 -2822
rect 117234 190894 117854 198000
rect 118374 197845 118434 199550
rect 120950 199550 121060 199610
rect 123448 199610 123508 200130
rect 125896 199610 125956 200130
rect 128480 199610 128540 200130
rect 130928 199610 130988 200130
rect 133512 199610 133572 200130
rect 123448 199550 123586 199610
rect 125896 199550 125978 199610
rect 128480 199550 128554 199610
rect 120950 198661 121010 199550
rect 123526 198661 123586 199550
rect 120947 198660 121013 198661
rect 120947 198596 120948 198660
rect 121012 198596 121013 198660
rect 120947 198595 121013 198596
rect 123523 198660 123589 198661
rect 123523 198596 123524 198660
rect 123588 198596 123589 198660
rect 123523 198595 123589 198596
rect 118371 197844 118437 197845
rect 118371 197780 118372 197844
rect 118436 197780 118437 197844
rect 118371 197779 118437 197780
rect 117234 190658 117266 190894
rect 117502 190658 117586 190894
rect 117822 190658 117854 190894
rect 117234 190574 117854 190658
rect 117234 190338 117266 190574
rect 117502 190338 117586 190574
rect 117822 190338 117854 190574
rect 117234 154894 117854 190338
rect 117234 154658 117266 154894
rect 117502 154658 117586 154894
rect 117822 154658 117854 154894
rect 117234 154574 117854 154658
rect 117234 154338 117266 154574
rect 117502 154338 117586 154574
rect 117822 154338 117854 154574
rect 117234 118894 117854 154338
rect 117234 118658 117266 118894
rect 117502 118658 117586 118894
rect 117822 118658 117854 118894
rect 117234 118574 117854 118658
rect 117234 118338 117266 118574
rect 117502 118338 117586 118574
rect 117822 118338 117854 118574
rect 117234 82894 117854 118338
rect 117234 82658 117266 82894
rect 117502 82658 117586 82894
rect 117822 82658 117854 82894
rect 117234 82574 117854 82658
rect 117234 82338 117266 82574
rect 117502 82338 117586 82574
rect 117822 82338 117854 82574
rect 117234 46894 117854 82338
rect 117234 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 117854 46894
rect 117234 46574 117854 46658
rect 117234 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 117854 46574
rect 117234 10894 117854 46338
rect 117234 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 117854 10894
rect 117234 10574 117854 10658
rect 117234 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 117854 10574
rect 117234 -4186 117854 10338
rect 117234 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 117854 -4186
rect 117234 -4506 117854 -4422
rect 117234 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 117854 -4506
rect 117234 -5734 117854 -4742
rect 120954 194614 121574 198000
rect 125918 197709 125978 199550
rect 128494 198661 128554 199550
rect 130886 199550 130988 199610
rect 133462 199550 133572 199610
rect 135960 199610 136020 200130
rect 138544 199610 138604 200130
rect 140992 199610 141052 200130
rect 143440 199610 143500 200130
rect 135960 199550 136098 199610
rect 138544 199550 138674 199610
rect 140992 199550 141066 199610
rect 130886 198661 130946 199550
rect 128491 198660 128557 198661
rect 128491 198596 128492 198660
rect 128556 198596 128557 198660
rect 128491 198595 128557 198596
rect 130883 198660 130949 198661
rect 130883 198596 130884 198660
rect 130948 198596 130949 198660
rect 130883 198595 130949 198596
rect 125915 197708 125981 197709
rect 125915 197644 125916 197708
rect 125980 197644 125981 197708
rect 125915 197643 125981 197644
rect 120954 194378 120986 194614
rect 121222 194378 121306 194614
rect 121542 194378 121574 194614
rect 120954 194294 121574 194378
rect 120954 194058 120986 194294
rect 121222 194058 121306 194294
rect 121542 194058 121574 194294
rect 120954 158614 121574 194058
rect 120954 158378 120986 158614
rect 121222 158378 121306 158614
rect 121542 158378 121574 158614
rect 120954 158294 121574 158378
rect 120954 158058 120986 158294
rect 121222 158058 121306 158294
rect 121542 158058 121574 158294
rect 120954 122614 121574 158058
rect 120954 122378 120986 122614
rect 121222 122378 121306 122614
rect 121542 122378 121574 122614
rect 120954 122294 121574 122378
rect 120954 122058 120986 122294
rect 121222 122058 121306 122294
rect 121542 122058 121574 122294
rect 120954 86614 121574 122058
rect 120954 86378 120986 86614
rect 121222 86378 121306 86614
rect 121542 86378 121574 86614
rect 120954 86294 121574 86378
rect 120954 86058 120986 86294
rect 121222 86058 121306 86294
rect 121542 86058 121574 86294
rect 120954 50614 121574 86058
rect 120954 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 121574 50614
rect 120954 50294 121574 50378
rect 120954 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 121574 50294
rect 120954 14614 121574 50058
rect 120954 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 121574 14614
rect 120954 14294 121574 14378
rect 120954 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 121574 14294
rect 102954 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 103574 -7066
rect 102954 -7386 103574 -7302
rect 102954 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 103574 -7386
rect 102954 -7654 103574 -7622
rect 120954 -6106 121574 14058
rect 127794 165454 128414 198000
rect 127794 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 128414 165454
rect 127794 165134 128414 165218
rect 127794 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 128414 165134
rect 127794 129454 128414 164898
rect 127794 129218 127826 129454
rect 128062 129218 128146 129454
rect 128382 129218 128414 129454
rect 127794 129134 128414 129218
rect 127794 128898 127826 129134
rect 128062 128898 128146 129134
rect 128382 128898 128414 129134
rect 127794 93454 128414 128898
rect 127794 93218 127826 93454
rect 128062 93218 128146 93454
rect 128382 93218 128414 93454
rect 127794 93134 128414 93218
rect 127794 92898 127826 93134
rect 128062 92898 128146 93134
rect 128382 92898 128414 93134
rect 127794 57454 128414 92898
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -1306 128414 20898
rect 127794 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 128414 -1306
rect 127794 -1626 128414 -1542
rect 127794 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 128414 -1626
rect 127794 -1894 128414 -1862
rect 131514 169174 132134 198000
rect 133462 197709 133522 199550
rect 136038 198661 136098 199550
rect 138614 198661 138674 199550
rect 136035 198660 136101 198661
rect 136035 198596 136036 198660
rect 136100 198596 136101 198660
rect 136035 198595 136101 198596
rect 138611 198660 138677 198661
rect 138611 198596 138612 198660
rect 138676 198596 138677 198660
rect 138611 198595 138677 198596
rect 133459 197708 133525 197709
rect 133459 197644 133460 197708
rect 133524 197644 133525 197708
rect 133459 197643 133525 197644
rect 131514 168938 131546 169174
rect 131782 168938 131866 169174
rect 132102 168938 132134 169174
rect 131514 168854 132134 168938
rect 131514 168618 131546 168854
rect 131782 168618 131866 168854
rect 132102 168618 132134 168854
rect 131514 133174 132134 168618
rect 131514 132938 131546 133174
rect 131782 132938 131866 133174
rect 132102 132938 132134 133174
rect 131514 132854 132134 132938
rect 131514 132618 131546 132854
rect 131782 132618 131866 132854
rect 132102 132618 132134 132854
rect 131514 97174 132134 132618
rect 131514 96938 131546 97174
rect 131782 96938 131866 97174
rect 132102 96938 132134 97174
rect 131514 96854 132134 96938
rect 131514 96618 131546 96854
rect 131782 96618 131866 96854
rect 132102 96618 132134 96854
rect 131514 61174 132134 96618
rect 131514 60938 131546 61174
rect 131782 60938 131866 61174
rect 132102 60938 132134 61174
rect 131514 60854 132134 60938
rect 131514 60618 131546 60854
rect 131782 60618 131866 60854
rect 132102 60618 132134 60854
rect 131514 25174 132134 60618
rect 131514 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 132134 25174
rect 131514 24854 132134 24938
rect 131514 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 132134 24854
rect 131514 -3226 132134 24618
rect 131514 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 132134 -3226
rect 131514 -3546 132134 -3462
rect 131514 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 132134 -3546
rect 131514 -3814 132134 -3782
rect 135234 172894 135854 198000
rect 135234 172658 135266 172894
rect 135502 172658 135586 172894
rect 135822 172658 135854 172894
rect 135234 172574 135854 172658
rect 135234 172338 135266 172574
rect 135502 172338 135586 172574
rect 135822 172338 135854 172574
rect 135234 136894 135854 172338
rect 135234 136658 135266 136894
rect 135502 136658 135586 136894
rect 135822 136658 135854 136894
rect 135234 136574 135854 136658
rect 135234 136338 135266 136574
rect 135502 136338 135586 136574
rect 135822 136338 135854 136574
rect 135234 100894 135854 136338
rect 135234 100658 135266 100894
rect 135502 100658 135586 100894
rect 135822 100658 135854 100894
rect 135234 100574 135854 100658
rect 135234 100338 135266 100574
rect 135502 100338 135586 100574
rect 135822 100338 135854 100574
rect 135234 64894 135854 100338
rect 135234 64658 135266 64894
rect 135502 64658 135586 64894
rect 135822 64658 135854 64894
rect 135234 64574 135854 64658
rect 135234 64338 135266 64574
rect 135502 64338 135586 64574
rect 135822 64338 135854 64574
rect 135234 28894 135854 64338
rect 135234 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 135854 28894
rect 135234 28574 135854 28658
rect 135234 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 135854 28574
rect 135234 -5146 135854 28338
rect 135234 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 135854 -5146
rect 135234 -5466 135854 -5382
rect 135234 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 135854 -5466
rect 135234 -5734 135854 -5702
rect 138954 176614 139574 198000
rect 141006 197981 141066 199550
rect 143398 199550 143500 199610
rect 145888 199610 145948 200130
rect 148472 199610 148532 200130
rect 150920 199610 150980 200130
rect 153368 199610 153428 200130
rect 155952 199610 156012 200130
rect 173224 199610 173284 200130
rect 145888 199550 146034 199610
rect 148472 199550 148610 199610
rect 150920 199550 151002 199610
rect 143398 198661 143458 199550
rect 145974 198661 146034 199550
rect 148550 198661 148610 199550
rect 150942 199477 151002 199550
rect 153334 199550 153428 199610
rect 155910 199550 156012 199610
rect 173206 199550 173284 199610
rect 173360 199610 173420 200130
rect 173360 199550 173450 199610
rect 150939 199476 151005 199477
rect 150939 199412 150940 199476
rect 151004 199412 151005 199476
rect 150939 199411 151005 199412
rect 153334 198661 153394 199550
rect 143395 198660 143461 198661
rect 143395 198596 143396 198660
rect 143460 198596 143461 198660
rect 143395 198595 143461 198596
rect 145971 198660 146037 198661
rect 145971 198596 145972 198660
rect 146036 198596 146037 198660
rect 145971 198595 146037 198596
rect 148547 198660 148613 198661
rect 148547 198596 148548 198660
rect 148612 198596 148613 198660
rect 148547 198595 148613 198596
rect 153331 198660 153397 198661
rect 153331 198596 153332 198660
rect 153396 198596 153397 198660
rect 153331 198595 153397 198596
rect 141003 197980 141069 197981
rect 141003 197916 141004 197980
rect 141068 197916 141069 197980
rect 141003 197915 141069 197916
rect 138954 176378 138986 176614
rect 139222 176378 139306 176614
rect 139542 176378 139574 176614
rect 138954 176294 139574 176378
rect 138954 176058 138986 176294
rect 139222 176058 139306 176294
rect 139542 176058 139574 176294
rect 138954 140614 139574 176058
rect 138954 140378 138986 140614
rect 139222 140378 139306 140614
rect 139542 140378 139574 140614
rect 138954 140294 139574 140378
rect 138954 140058 138986 140294
rect 139222 140058 139306 140294
rect 139542 140058 139574 140294
rect 138954 104614 139574 140058
rect 138954 104378 138986 104614
rect 139222 104378 139306 104614
rect 139542 104378 139574 104614
rect 138954 104294 139574 104378
rect 138954 104058 138986 104294
rect 139222 104058 139306 104294
rect 139542 104058 139574 104294
rect 138954 68614 139574 104058
rect 138954 68378 138986 68614
rect 139222 68378 139306 68614
rect 139542 68378 139574 68614
rect 138954 68294 139574 68378
rect 138954 68058 138986 68294
rect 139222 68058 139306 68294
rect 139542 68058 139574 68294
rect 138954 32614 139574 68058
rect 138954 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 139574 32614
rect 138954 32294 139574 32378
rect 138954 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 139574 32294
rect 120954 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 121574 -6106
rect 120954 -6426 121574 -6342
rect 120954 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 121574 -6426
rect 120954 -7654 121574 -6662
rect 138954 -7066 139574 32058
rect 145794 183454 146414 198000
rect 145794 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 146414 183454
rect 145794 183134 146414 183218
rect 145794 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 146414 183134
rect 145794 147454 146414 182898
rect 145794 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 146414 147454
rect 145794 147134 146414 147218
rect 145794 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 146414 147134
rect 145794 111454 146414 146898
rect 145794 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 146414 111454
rect 145794 111134 146414 111218
rect 145794 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 146414 111134
rect 145794 75454 146414 110898
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 145794 39454 146414 74898
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -1894 146414 -902
rect 149514 187174 150134 198000
rect 149514 186938 149546 187174
rect 149782 186938 149866 187174
rect 150102 186938 150134 187174
rect 149514 186854 150134 186938
rect 149514 186618 149546 186854
rect 149782 186618 149866 186854
rect 150102 186618 150134 186854
rect 149514 151174 150134 186618
rect 149514 150938 149546 151174
rect 149782 150938 149866 151174
rect 150102 150938 150134 151174
rect 149514 150854 150134 150938
rect 149514 150618 149546 150854
rect 149782 150618 149866 150854
rect 150102 150618 150134 150854
rect 149514 115174 150134 150618
rect 149514 114938 149546 115174
rect 149782 114938 149866 115174
rect 150102 114938 150134 115174
rect 149514 114854 150134 114938
rect 149514 114618 149546 114854
rect 149782 114618 149866 114854
rect 150102 114618 150134 114854
rect 149514 79174 150134 114618
rect 149514 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 150134 79174
rect 149514 78854 150134 78938
rect 149514 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 150134 78854
rect 149514 43174 150134 78618
rect 149514 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 150134 43174
rect 149514 42854 150134 42938
rect 149514 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 150134 42854
rect 149514 7174 150134 42618
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -2266 150134 6618
rect 149514 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 150134 -2266
rect 149514 -2586 150134 -2502
rect 149514 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 150134 -2586
rect 149514 -3814 150134 -2822
rect 153234 190894 153854 198000
rect 155910 197845 155970 199550
rect 155907 197844 155973 197845
rect 155907 197780 155908 197844
rect 155972 197780 155973 197844
rect 155907 197779 155973 197780
rect 153234 190658 153266 190894
rect 153502 190658 153586 190894
rect 153822 190658 153854 190894
rect 153234 190574 153854 190658
rect 153234 190338 153266 190574
rect 153502 190338 153586 190574
rect 153822 190338 153854 190574
rect 153234 154894 153854 190338
rect 153234 154658 153266 154894
rect 153502 154658 153586 154894
rect 153822 154658 153854 154894
rect 153234 154574 153854 154658
rect 153234 154338 153266 154574
rect 153502 154338 153586 154574
rect 153822 154338 153854 154574
rect 153234 118894 153854 154338
rect 153234 118658 153266 118894
rect 153502 118658 153586 118894
rect 153822 118658 153854 118894
rect 153234 118574 153854 118658
rect 153234 118338 153266 118574
rect 153502 118338 153586 118574
rect 153822 118338 153854 118574
rect 153234 82894 153854 118338
rect 153234 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 153854 82894
rect 153234 82574 153854 82658
rect 153234 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 153854 82574
rect 153234 46894 153854 82338
rect 153234 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 153854 46894
rect 153234 46574 153854 46658
rect 153234 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 153854 46574
rect 153234 10894 153854 46338
rect 153234 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 153854 10894
rect 153234 10574 153854 10658
rect 153234 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 153854 10574
rect 153234 -4186 153854 10338
rect 153234 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 153854 -4186
rect 153234 -4506 153854 -4422
rect 153234 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 153854 -4506
rect 153234 -5734 153854 -4742
rect 156954 194614 157574 198000
rect 156954 194378 156986 194614
rect 157222 194378 157306 194614
rect 157542 194378 157574 194614
rect 156954 194294 157574 194378
rect 156954 194058 156986 194294
rect 157222 194058 157306 194294
rect 157542 194058 157574 194294
rect 156954 158614 157574 194058
rect 156954 158378 156986 158614
rect 157222 158378 157306 158614
rect 157542 158378 157574 158614
rect 156954 158294 157574 158378
rect 156954 158058 156986 158294
rect 157222 158058 157306 158294
rect 157542 158058 157574 158294
rect 156954 122614 157574 158058
rect 156954 122378 156986 122614
rect 157222 122378 157306 122614
rect 157542 122378 157574 122614
rect 156954 122294 157574 122378
rect 156954 122058 156986 122294
rect 157222 122058 157306 122294
rect 157542 122058 157574 122294
rect 156954 86614 157574 122058
rect 156954 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 157574 86614
rect 156954 86294 157574 86378
rect 156954 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 157574 86294
rect 156954 50614 157574 86058
rect 156954 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 157574 50614
rect 156954 50294 157574 50378
rect 156954 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 157574 50294
rect 156954 14614 157574 50058
rect 156954 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 157574 14614
rect 156954 14294 157574 14378
rect 156954 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 157574 14294
rect 138954 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 139574 -7066
rect 138954 -7386 139574 -7302
rect 138954 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 139574 -7386
rect 138954 -7654 139574 -7622
rect 156954 -6106 157574 14058
rect 163794 165454 164414 198000
rect 163794 165218 163826 165454
rect 164062 165218 164146 165454
rect 164382 165218 164414 165454
rect 163794 165134 164414 165218
rect 163794 164898 163826 165134
rect 164062 164898 164146 165134
rect 164382 164898 164414 165134
rect 163794 129454 164414 164898
rect 163794 129218 163826 129454
rect 164062 129218 164146 129454
rect 164382 129218 164414 129454
rect 163794 129134 164414 129218
rect 163794 128898 163826 129134
rect 164062 128898 164146 129134
rect 164382 128898 164414 129134
rect 163794 93454 164414 128898
rect 163794 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 164414 93454
rect 163794 93134 164414 93218
rect 163794 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 164414 93134
rect 163794 57454 164414 92898
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -1306 164414 20898
rect 163794 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 164414 -1306
rect 163794 -1626 164414 -1542
rect 163794 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 164414 -1626
rect 163794 -1894 164414 -1862
rect 167514 169174 168134 198000
rect 167514 168938 167546 169174
rect 167782 168938 167866 169174
rect 168102 168938 168134 169174
rect 167514 168854 168134 168938
rect 167514 168618 167546 168854
rect 167782 168618 167866 168854
rect 168102 168618 168134 168854
rect 167514 133174 168134 168618
rect 167514 132938 167546 133174
rect 167782 132938 167866 133174
rect 168102 132938 168134 133174
rect 167514 132854 168134 132938
rect 167514 132618 167546 132854
rect 167782 132618 167866 132854
rect 168102 132618 168134 132854
rect 167514 97174 168134 132618
rect 167514 96938 167546 97174
rect 167782 96938 167866 97174
rect 168102 96938 168134 97174
rect 167514 96854 168134 96938
rect 167514 96618 167546 96854
rect 167782 96618 167866 96854
rect 168102 96618 168134 96854
rect 167514 61174 168134 96618
rect 167514 60938 167546 61174
rect 167782 60938 167866 61174
rect 168102 60938 168134 61174
rect 167514 60854 168134 60938
rect 167514 60618 167546 60854
rect 167782 60618 167866 60854
rect 168102 60618 168134 60854
rect 167514 25174 168134 60618
rect 167514 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 168134 25174
rect 167514 24854 168134 24938
rect 167514 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 168134 24854
rect 167514 -3226 168134 24618
rect 167514 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 168134 -3226
rect 167514 -3546 168134 -3462
rect 167514 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 168134 -3546
rect 167514 -3814 168134 -3782
rect 171234 172894 171854 198000
rect 173206 197845 173266 199550
rect 173390 198661 173450 199550
rect 186822 198933 186882 277475
rect 187003 271964 187069 271965
rect 187003 271900 187004 271964
rect 187068 271900 187069 271964
rect 187003 271899 187069 271900
rect 186819 198932 186885 198933
rect 186819 198868 186820 198932
rect 186884 198868 186885 198932
rect 186819 198867 186885 198868
rect 173387 198660 173453 198661
rect 173387 198596 173388 198660
rect 173452 198596 173453 198660
rect 173387 198595 173453 198596
rect 187006 198253 187066 271899
rect 187190 255373 187250 285907
rect 188291 279036 188357 279037
rect 188291 278972 188292 279036
rect 188356 278972 188357 279036
rect 188291 278971 188357 278972
rect 187187 255372 187253 255373
rect 187187 255308 187188 255372
rect 187252 255308 187253 255372
rect 187187 255307 187253 255308
rect 187187 205732 187253 205733
rect 187187 205668 187188 205732
rect 187252 205668 187253 205732
rect 187187 205667 187253 205668
rect 187003 198252 187069 198253
rect 187003 198188 187004 198252
rect 187068 198188 187069 198252
rect 187003 198187 187069 198188
rect 187190 198117 187250 205667
rect 187187 198116 187253 198117
rect 187187 198052 187188 198116
rect 187252 198052 187253 198116
rect 187187 198051 187253 198052
rect 173203 197844 173269 197845
rect 173203 197780 173204 197844
rect 173268 197780 173269 197844
rect 173203 197779 173269 197780
rect 171234 172658 171266 172894
rect 171502 172658 171586 172894
rect 171822 172658 171854 172894
rect 171234 172574 171854 172658
rect 171234 172338 171266 172574
rect 171502 172338 171586 172574
rect 171822 172338 171854 172574
rect 171234 136894 171854 172338
rect 171234 136658 171266 136894
rect 171502 136658 171586 136894
rect 171822 136658 171854 136894
rect 171234 136574 171854 136658
rect 171234 136338 171266 136574
rect 171502 136338 171586 136574
rect 171822 136338 171854 136574
rect 171234 100894 171854 136338
rect 171234 100658 171266 100894
rect 171502 100658 171586 100894
rect 171822 100658 171854 100894
rect 171234 100574 171854 100658
rect 171234 100338 171266 100574
rect 171502 100338 171586 100574
rect 171822 100338 171854 100574
rect 171234 64894 171854 100338
rect 171234 64658 171266 64894
rect 171502 64658 171586 64894
rect 171822 64658 171854 64894
rect 171234 64574 171854 64658
rect 171234 64338 171266 64574
rect 171502 64338 171586 64574
rect 171822 64338 171854 64574
rect 171234 28894 171854 64338
rect 171234 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 171854 28894
rect 171234 28574 171854 28658
rect 171234 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 171854 28574
rect 171234 -5146 171854 28338
rect 171234 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 171854 -5146
rect 171234 -5466 171854 -5382
rect 171234 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 171854 -5466
rect 171234 -5734 171854 -5702
rect 174954 176614 175574 198000
rect 174954 176378 174986 176614
rect 175222 176378 175306 176614
rect 175542 176378 175574 176614
rect 174954 176294 175574 176378
rect 174954 176058 174986 176294
rect 175222 176058 175306 176294
rect 175542 176058 175574 176294
rect 174954 140614 175574 176058
rect 174954 140378 174986 140614
rect 175222 140378 175306 140614
rect 175542 140378 175574 140614
rect 174954 140294 175574 140378
rect 174954 140058 174986 140294
rect 175222 140058 175306 140294
rect 175542 140058 175574 140294
rect 174954 104614 175574 140058
rect 174954 104378 174986 104614
rect 175222 104378 175306 104614
rect 175542 104378 175574 104614
rect 174954 104294 175574 104378
rect 174954 104058 174986 104294
rect 175222 104058 175306 104294
rect 175542 104058 175574 104294
rect 174954 68614 175574 104058
rect 174954 68378 174986 68614
rect 175222 68378 175306 68614
rect 175542 68378 175574 68614
rect 174954 68294 175574 68378
rect 174954 68058 174986 68294
rect 175222 68058 175306 68294
rect 175542 68058 175574 68294
rect 174954 32614 175574 68058
rect 174954 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 175574 32614
rect 174954 32294 175574 32378
rect 174954 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 175574 32294
rect 156954 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 157574 -6106
rect 156954 -6426 157574 -6342
rect 156954 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 157574 -6426
rect 156954 -7654 157574 -6662
rect 174954 -7066 175574 32058
rect 181794 183454 182414 198000
rect 181794 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 182414 183454
rect 181794 183134 182414 183218
rect 181794 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 182414 183134
rect 181794 147454 182414 182898
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 111454 182414 146898
rect 181794 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 182414 111454
rect 181794 111134 182414 111218
rect 181794 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 182414 111134
rect 181794 75454 182414 110898
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 181794 39454 182414 74898
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -1894 182414 -902
rect 185514 187174 186134 198000
rect 188294 196757 188354 278971
rect 188475 276180 188541 276181
rect 188475 276116 188476 276180
rect 188540 276116 188541 276180
rect 188475 276115 188541 276116
rect 188478 197981 188538 276115
rect 188659 273460 188725 273461
rect 188659 273396 188660 273460
rect 188724 273396 188725 273460
rect 188659 273395 188725 273396
rect 188475 197980 188541 197981
rect 188475 197916 188476 197980
rect 188540 197916 188541 197980
rect 188475 197915 188541 197916
rect 188662 196893 188722 273395
rect 189234 262894 189854 298338
rect 189234 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 189854 262894
rect 189234 262574 189854 262658
rect 189234 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 189854 262574
rect 189234 226894 189854 262338
rect 189234 226658 189266 226894
rect 189502 226658 189586 226894
rect 189822 226658 189854 226894
rect 189234 226574 189854 226658
rect 189234 226338 189266 226574
rect 189502 226338 189586 226574
rect 189822 226338 189854 226574
rect 188659 196892 188725 196893
rect 188659 196828 188660 196892
rect 188724 196828 188725 196892
rect 188659 196827 188725 196828
rect 188291 196756 188357 196757
rect 188291 196692 188292 196756
rect 188356 196692 188357 196756
rect 188291 196691 188357 196692
rect 185514 186938 185546 187174
rect 185782 186938 185866 187174
rect 186102 186938 186134 187174
rect 185514 186854 186134 186938
rect 185514 186618 185546 186854
rect 185782 186618 185866 186854
rect 186102 186618 186134 186854
rect 185514 151174 186134 186618
rect 185514 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 186134 151174
rect 185514 150854 186134 150938
rect 185514 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 186134 150854
rect 185514 115174 186134 150618
rect 185514 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 186134 115174
rect 185514 114854 186134 114938
rect 185514 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 186134 114854
rect 185514 79174 186134 114618
rect 185514 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 186134 79174
rect 185514 78854 186134 78938
rect 185514 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 186134 78854
rect 185514 43174 186134 78618
rect 185514 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 186134 43174
rect 185514 42854 186134 42938
rect 185514 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 186134 42854
rect 185514 7174 186134 42618
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 185514 -2266 186134 6618
rect 185514 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 186134 -2266
rect 185514 -2586 186134 -2502
rect 185514 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 186134 -2586
rect 185514 -3814 186134 -2822
rect 189234 190894 189854 226338
rect 189234 190658 189266 190894
rect 189502 190658 189586 190894
rect 189822 190658 189854 190894
rect 189234 190574 189854 190658
rect 189234 190338 189266 190574
rect 189502 190338 189586 190574
rect 189822 190338 189854 190574
rect 189234 154894 189854 190338
rect 189234 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 189854 154894
rect 189234 154574 189854 154658
rect 189234 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 189854 154574
rect 189234 118894 189854 154338
rect 189234 118658 189266 118894
rect 189502 118658 189586 118894
rect 189822 118658 189854 118894
rect 189234 118574 189854 118658
rect 189234 118338 189266 118574
rect 189502 118338 189586 118574
rect 189822 118338 189854 118574
rect 189234 82894 189854 118338
rect 189234 82658 189266 82894
rect 189502 82658 189586 82894
rect 189822 82658 189854 82894
rect 189234 82574 189854 82658
rect 189234 82338 189266 82574
rect 189502 82338 189586 82574
rect 189822 82338 189854 82574
rect 189234 46894 189854 82338
rect 189234 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 189854 46894
rect 189234 46574 189854 46658
rect 189234 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 189854 46574
rect 189234 10894 189854 46338
rect 189234 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 189854 10894
rect 189234 10574 189854 10658
rect 189234 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 189854 10574
rect 189234 -4186 189854 10338
rect 189234 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 189854 -4186
rect 189234 -4506 189854 -4422
rect 189234 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 189854 -4506
rect 189234 -5734 189854 -4742
rect 192954 698614 193574 710042
rect 210954 711558 211574 711590
rect 210954 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 211574 711558
rect 210954 711238 211574 711322
rect 210954 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 211574 711238
rect 207234 709638 207854 709670
rect 207234 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 207854 709638
rect 207234 709318 207854 709402
rect 207234 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 207854 709318
rect 203514 707718 204134 707750
rect 203514 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 204134 707718
rect 203514 707398 204134 707482
rect 203514 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 204134 707398
rect 192954 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 193574 698614
rect 192954 698294 193574 698378
rect 192954 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 193574 698294
rect 192954 662614 193574 698058
rect 192954 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 193574 662614
rect 192954 662294 193574 662378
rect 192954 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 193574 662294
rect 192954 626614 193574 662058
rect 192954 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 193574 626614
rect 192954 626294 193574 626378
rect 192954 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 193574 626294
rect 192954 590614 193574 626058
rect 192954 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 193574 590614
rect 192954 590294 193574 590378
rect 192954 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 193574 590294
rect 192954 554614 193574 590058
rect 192954 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 193574 554614
rect 192954 554294 193574 554378
rect 192954 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 193574 554294
rect 192954 518614 193574 554058
rect 192954 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 193574 518614
rect 192954 518294 193574 518378
rect 192954 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 193574 518294
rect 192954 482614 193574 518058
rect 192954 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 193574 482614
rect 192954 482294 193574 482378
rect 192954 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 193574 482294
rect 192954 446614 193574 482058
rect 192954 446378 192986 446614
rect 193222 446378 193306 446614
rect 193542 446378 193574 446614
rect 192954 446294 193574 446378
rect 192954 446058 192986 446294
rect 193222 446058 193306 446294
rect 193542 446058 193574 446294
rect 192954 410614 193574 446058
rect 192954 410378 192986 410614
rect 193222 410378 193306 410614
rect 193542 410378 193574 410614
rect 192954 410294 193574 410378
rect 192954 410058 192986 410294
rect 193222 410058 193306 410294
rect 193542 410058 193574 410294
rect 192954 374614 193574 410058
rect 192954 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 193574 374614
rect 192954 374294 193574 374378
rect 192954 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 193574 374294
rect 192954 338614 193574 374058
rect 192954 338378 192986 338614
rect 193222 338378 193306 338614
rect 193542 338378 193574 338614
rect 192954 338294 193574 338378
rect 192954 338058 192986 338294
rect 193222 338058 193306 338294
rect 193542 338058 193574 338294
rect 192954 302614 193574 338058
rect 192954 302378 192986 302614
rect 193222 302378 193306 302614
rect 193542 302378 193574 302614
rect 192954 302294 193574 302378
rect 192954 302058 192986 302294
rect 193222 302058 193306 302294
rect 193542 302058 193574 302294
rect 192954 266614 193574 302058
rect 192954 266378 192986 266614
rect 193222 266378 193306 266614
rect 193542 266378 193574 266614
rect 192954 266294 193574 266378
rect 192954 266058 192986 266294
rect 193222 266058 193306 266294
rect 193542 266058 193574 266294
rect 192954 230614 193574 266058
rect 192954 230378 192986 230614
rect 193222 230378 193306 230614
rect 193542 230378 193574 230614
rect 192954 230294 193574 230378
rect 192954 230058 192986 230294
rect 193222 230058 193306 230294
rect 193542 230058 193574 230294
rect 192954 194614 193574 230058
rect 192954 194378 192986 194614
rect 193222 194378 193306 194614
rect 193542 194378 193574 194614
rect 192954 194294 193574 194378
rect 192954 194058 192986 194294
rect 193222 194058 193306 194294
rect 193542 194058 193574 194294
rect 192954 158614 193574 194058
rect 192954 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 193574 158614
rect 192954 158294 193574 158378
rect 192954 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 193574 158294
rect 192954 122614 193574 158058
rect 192954 122378 192986 122614
rect 193222 122378 193306 122614
rect 193542 122378 193574 122614
rect 192954 122294 193574 122378
rect 192954 122058 192986 122294
rect 193222 122058 193306 122294
rect 193542 122058 193574 122294
rect 192954 86614 193574 122058
rect 192954 86378 192986 86614
rect 193222 86378 193306 86614
rect 193542 86378 193574 86614
rect 192954 86294 193574 86378
rect 192954 86058 192986 86294
rect 193222 86058 193306 86294
rect 193542 86058 193574 86294
rect 192954 50614 193574 86058
rect 192954 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 193574 50614
rect 192954 50294 193574 50378
rect 192954 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 193574 50294
rect 192954 14614 193574 50058
rect 192954 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 193574 14614
rect 192954 14294 193574 14378
rect 192954 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 193574 14294
rect 174954 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 175574 -7066
rect 174954 -7386 175574 -7302
rect 174954 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 175574 -7386
rect 174954 -7654 175574 -7622
rect 192954 -6106 193574 14058
rect 199794 705798 200414 705830
rect 199794 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 200414 705798
rect 199794 705478 200414 705562
rect 199794 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 200414 705478
rect 199794 669454 200414 705242
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 561454 200414 596898
rect 199794 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 200414 561454
rect 199794 561134 200414 561218
rect 199794 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 200414 561134
rect 199794 525454 200414 560898
rect 199794 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 200414 525454
rect 199794 525134 200414 525218
rect 199794 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 200414 525134
rect 199794 489454 200414 524898
rect 199794 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 200414 489454
rect 199794 489134 200414 489218
rect 199794 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 200414 489134
rect 199794 453454 200414 488898
rect 199794 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 200414 453454
rect 199794 453134 200414 453218
rect 199794 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 200414 453134
rect 199794 417454 200414 452898
rect 199794 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 200414 417454
rect 199794 417134 200414 417218
rect 199794 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 200414 417134
rect 199794 381454 200414 416898
rect 199794 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 200414 381454
rect 199794 381134 200414 381218
rect 199794 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 200414 381134
rect 199794 345454 200414 380898
rect 199794 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 200414 345454
rect 199794 345134 200414 345218
rect 199794 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 200414 345134
rect 199794 309454 200414 344898
rect 199794 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 200414 309454
rect 199794 309134 200414 309218
rect 199794 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 200414 309134
rect 199794 273454 200414 308898
rect 199794 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 200414 273454
rect 199794 273134 200414 273218
rect 199794 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 200414 273134
rect 199794 237454 200414 272898
rect 199794 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 200414 237454
rect 199794 237134 200414 237218
rect 199794 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 200414 237134
rect 199794 201454 200414 236898
rect 199794 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 200414 201454
rect 199794 201134 200414 201218
rect 199794 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 200414 201134
rect 199794 165454 200414 200898
rect 199794 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 200414 165454
rect 199794 165134 200414 165218
rect 199794 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 200414 165134
rect 199794 129454 200414 164898
rect 199794 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 200414 129454
rect 199794 129134 200414 129218
rect 199794 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 200414 129134
rect 199794 93454 200414 128898
rect 199794 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 200414 93454
rect 199794 93134 200414 93218
rect 199794 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 200414 93134
rect 199794 57454 200414 92898
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -1306 200414 20898
rect 199794 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 200414 -1306
rect 199794 -1626 200414 -1542
rect 199794 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 200414 -1626
rect 199794 -1894 200414 -1862
rect 203514 673174 204134 707162
rect 203514 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 204134 673174
rect 203514 672854 204134 672938
rect 203514 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 204134 672854
rect 203514 637174 204134 672618
rect 203514 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 204134 637174
rect 203514 636854 204134 636938
rect 203514 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 204134 636854
rect 203514 601174 204134 636618
rect 203514 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 204134 601174
rect 203514 600854 204134 600938
rect 203514 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 204134 600854
rect 203514 565174 204134 600618
rect 203514 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 204134 565174
rect 203514 564854 204134 564938
rect 203514 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 204134 564854
rect 203514 529174 204134 564618
rect 203514 528938 203546 529174
rect 203782 528938 203866 529174
rect 204102 528938 204134 529174
rect 203514 528854 204134 528938
rect 203514 528618 203546 528854
rect 203782 528618 203866 528854
rect 204102 528618 204134 528854
rect 203514 493174 204134 528618
rect 203514 492938 203546 493174
rect 203782 492938 203866 493174
rect 204102 492938 204134 493174
rect 203514 492854 204134 492938
rect 203514 492618 203546 492854
rect 203782 492618 203866 492854
rect 204102 492618 204134 492854
rect 203514 457174 204134 492618
rect 203514 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 204134 457174
rect 203514 456854 204134 456938
rect 203514 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 204134 456854
rect 203514 421174 204134 456618
rect 203514 420938 203546 421174
rect 203782 420938 203866 421174
rect 204102 420938 204134 421174
rect 203514 420854 204134 420938
rect 203514 420618 203546 420854
rect 203782 420618 203866 420854
rect 204102 420618 204134 420854
rect 203514 385174 204134 420618
rect 203514 384938 203546 385174
rect 203782 384938 203866 385174
rect 204102 384938 204134 385174
rect 203514 384854 204134 384938
rect 203514 384618 203546 384854
rect 203782 384618 203866 384854
rect 204102 384618 204134 384854
rect 203514 349174 204134 384618
rect 203514 348938 203546 349174
rect 203782 348938 203866 349174
rect 204102 348938 204134 349174
rect 203514 348854 204134 348938
rect 203514 348618 203546 348854
rect 203782 348618 203866 348854
rect 204102 348618 204134 348854
rect 203514 313174 204134 348618
rect 203514 312938 203546 313174
rect 203782 312938 203866 313174
rect 204102 312938 204134 313174
rect 203514 312854 204134 312938
rect 203514 312618 203546 312854
rect 203782 312618 203866 312854
rect 204102 312618 204134 312854
rect 203514 277174 204134 312618
rect 203514 276938 203546 277174
rect 203782 276938 203866 277174
rect 204102 276938 204134 277174
rect 203514 276854 204134 276938
rect 203514 276618 203546 276854
rect 203782 276618 203866 276854
rect 204102 276618 204134 276854
rect 203514 241174 204134 276618
rect 203514 240938 203546 241174
rect 203782 240938 203866 241174
rect 204102 240938 204134 241174
rect 203514 240854 204134 240938
rect 203514 240618 203546 240854
rect 203782 240618 203866 240854
rect 204102 240618 204134 240854
rect 203514 205174 204134 240618
rect 203514 204938 203546 205174
rect 203782 204938 203866 205174
rect 204102 204938 204134 205174
rect 203514 204854 204134 204938
rect 203514 204618 203546 204854
rect 203782 204618 203866 204854
rect 204102 204618 204134 204854
rect 203514 169174 204134 204618
rect 203514 168938 203546 169174
rect 203782 168938 203866 169174
rect 204102 168938 204134 169174
rect 203514 168854 204134 168938
rect 203514 168618 203546 168854
rect 203782 168618 203866 168854
rect 204102 168618 204134 168854
rect 203514 133174 204134 168618
rect 203514 132938 203546 133174
rect 203782 132938 203866 133174
rect 204102 132938 204134 133174
rect 203514 132854 204134 132938
rect 203514 132618 203546 132854
rect 203782 132618 203866 132854
rect 204102 132618 204134 132854
rect 203514 97174 204134 132618
rect 203514 96938 203546 97174
rect 203782 96938 203866 97174
rect 204102 96938 204134 97174
rect 203514 96854 204134 96938
rect 203514 96618 203546 96854
rect 203782 96618 203866 96854
rect 204102 96618 204134 96854
rect 203514 61174 204134 96618
rect 203514 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 204134 61174
rect 203514 60854 204134 60938
rect 203514 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 204134 60854
rect 203514 25174 204134 60618
rect 203514 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 204134 25174
rect 203514 24854 204134 24938
rect 203514 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 204134 24854
rect 203514 -3226 204134 24618
rect 203514 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 204134 -3226
rect 203514 -3546 204134 -3462
rect 203514 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 204134 -3546
rect 203514 -3814 204134 -3782
rect 207234 676894 207854 709082
rect 207234 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 207854 676894
rect 207234 676574 207854 676658
rect 207234 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 207854 676574
rect 207234 640894 207854 676338
rect 207234 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 207854 640894
rect 207234 640574 207854 640658
rect 207234 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 207854 640574
rect 207234 604894 207854 640338
rect 207234 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 207854 604894
rect 207234 604574 207854 604658
rect 207234 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 207854 604574
rect 207234 568894 207854 604338
rect 207234 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 207854 568894
rect 207234 568574 207854 568658
rect 207234 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 207854 568574
rect 207234 532894 207854 568338
rect 207234 532658 207266 532894
rect 207502 532658 207586 532894
rect 207822 532658 207854 532894
rect 207234 532574 207854 532658
rect 207234 532338 207266 532574
rect 207502 532338 207586 532574
rect 207822 532338 207854 532574
rect 207234 496894 207854 532338
rect 207234 496658 207266 496894
rect 207502 496658 207586 496894
rect 207822 496658 207854 496894
rect 207234 496574 207854 496658
rect 207234 496338 207266 496574
rect 207502 496338 207586 496574
rect 207822 496338 207854 496574
rect 207234 460894 207854 496338
rect 207234 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 207854 460894
rect 207234 460574 207854 460658
rect 207234 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 207854 460574
rect 207234 424894 207854 460338
rect 207234 424658 207266 424894
rect 207502 424658 207586 424894
rect 207822 424658 207854 424894
rect 207234 424574 207854 424658
rect 207234 424338 207266 424574
rect 207502 424338 207586 424574
rect 207822 424338 207854 424574
rect 207234 388894 207854 424338
rect 207234 388658 207266 388894
rect 207502 388658 207586 388894
rect 207822 388658 207854 388894
rect 207234 388574 207854 388658
rect 207234 388338 207266 388574
rect 207502 388338 207586 388574
rect 207822 388338 207854 388574
rect 207234 352894 207854 388338
rect 207234 352658 207266 352894
rect 207502 352658 207586 352894
rect 207822 352658 207854 352894
rect 207234 352574 207854 352658
rect 207234 352338 207266 352574
rect 207502 352338 207586 352574
rect 207822 352338 207854 352574
rect 207234 316894 207854 352338
rect 207234 316658 207266 316894
rect 207502 316658 207586 316894
rect 207822 316658 207854 316894
rect 207234 316574 207854 316658
rect 207234 316338 207266 316574
rect 207502 316338 207586 316574
rect 207822 316338 207854 316574
rect 207234 280894 207854 316338
rect 207234 280658 207266 280894
rect 207502 280658 207586 280894
rect 207822 280658 207854 280894
rect 207234 280574 207854 280658
rect 207234 280338 207266 280574
rect 207502 280338 207586 280574
rect 207822 280338 207854 280574
rect 207234 244894 207854 280338
rect 207234 244658 207266 244894
rect 207502 244658 207586 244894
rect 207822 244658 207854 244894
rect 207234 244574 207854 244658
rect 207234 244338 207266 244574
rect 207502 244338 207586 244574
rect 207822 244338 207854 244574
rect 207234 208894 207854 244338
rect 207234 208658 207266 208894
rect 207502 208658 207586 208894
rect 207822 208658 207854 208894
rect 207234 208574 207854 208658
rect 207234 208338 207266 208574
rect 207502 208338 207586 208574
rect 207822 208338 207854 208574
rect 207234 172894 207854 208338
rect 207234 172658 207266 172894
rect 207502 172658 207586 172894
rect 207822 172658 207854 172894
rect 207234 172574 207854 172658
rect 207234 172338 207266 172574
rect 207502 172338 207586 172574
rect 207822 172338 207854 172574
rect 207234 136894 207854 172338
rect 207234 136658 207266 136894
rect 207502 136658 207586 136894
rect 207822 136658 207854 136894
rect 207234 136574 207854 136658
rect 207234 136338 207266 136574
rect 207502 136338 207586 136574
rect 207822 136338 207854 136574
rect 207234 100894 207854 136338
rect 207234 100658 207266 100894
rect 207502 100658 207586 100894
rect 207822 100658 207854 100894
rect 207234 100574 207854 100658
rect 207234 100338 207266 100574
rect 207502 100338 207586 100574
rect 207822 100338 207854 100574
rect 207234 64894 207854 100338
rect 207234 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 207854 64894
rect 207234 64574 207854 64658
rect 207234 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 207854 64574
rect 207234 28894 207854 64338
rect 207234 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 207854 28894
rect 207234 28574 207854 28658
rect 207234 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 207854 28574
rect 207234 -5146 207854 28338
rect 207234 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 207854 -5146
rect 207234 -5466 207854 -5382
rect 207234 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 207854 -5466
rect 207234 -5734 207854 -5702
rect 210954 680614 211574 711002
rect 228954 710598 229574 711590
rect 228954 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 229574 710598
rect 228954 710278 229574 710362
rect 228954 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 229574 710278
rect 225234 708678 225854 709670
rect 225234 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 225854 708678
rect 225234 708358 225854 708442
rect 225234 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 225854 708358
rect 221514 706758 222134 707750
rect 221514 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 222134 706758
rect 221514 706438 222134 706522
rect 221514 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 222134 706438
rect 210954 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 211574 680614
rect 210954 680294 211574 680378
rect 210954 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 211574 680294
rect 210954 644614 211574 680058
rect 210954 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 211574 644614
rect 210954 644294 211574 644378
rect 210954 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 211574 644294
rect 210954 608614 211574 644058
rect 210954 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 211574 608614
rect 210954 608294 211574 608378
rect 210954 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 211574 608294
rect 210954 572614 211574 608058
rect 210954 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 211574 572614
rect 210954 572294 211574 572378
rect 210954 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 211574 572294
rect 210954 536614 211574 572058
rect 210954 536378 210986 536614
rect 211222 536378 211306 536614
rect 211542 536378 211574 536614
rect 210954 536294 211574 536378
rect 210954 536058 210986 536294
rect 211222 536058 211306 536294
rect 211542 536058 211574 536294
rect 210954 500614 211574 536058
rect 210954 500378 210986 500614
rect 211222 500378 211306 500614
rect 211542 500378 211574 500614
rect 210954 500294 211574 500378
rect 210954 500058 210986 500294
rect 211222 500058 211306 500294
rect 211542 500058 211574 500294
rect 210954 464614 211574 500058
rect 210954 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 211574 464614
rect 210954 464294 211574 464378
rect 210954 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 211574 464294
rect 210954 428614 211574 464058
rect 210954 428378 210986 428614
rect 211222 428378 211306 428614
rect 211542 428378 211574 428614
rect 210954 428294 211574 428378
rect 210954 428058 210986 428294
rect 211222 428058 211306 428294
rect 211542 428058 211574 428294
rect 210954 392614 211574 428058
rect 210954 392378 210986 392614
rect 211222 392378 211306 392614
rect 211542 392378 211574 392614
rect 210954 392294 211574 392378
rect 210954 392058 210986 392294
rect 211222 392058 211306 392294
rect 211542 392058 211574 392294
rect 210954 356614 211574 392058
rect 210954 356378 210986 356614
rect 211222 356378 211306 356614
rect 211542 356378 211574 356614
rect 210954 356294 211574 356378
rect 210954 356058 210986 356294
rect 211222 356058 211306 356294
rect 211542 356058 211574 356294
rect 210954 320614 211574 356058
rect 210954 320378 210986 320614
rect 211222 320378 211306 320614
rect 211542 320378 211574 320614
rect 210954 320294 211574 320378
rect 210954 320058 210986 320294
rect 211222 320058 211306 320294
rect 211542 320058 211574 320294
rect 210954 284614 211574 320058
rect 210954 284378 210986 284614
rect 211222 284378 211306 284614
rect 211542 284378 211574 284614
rect 210954 284294 211574 284378
rect 210954 284058 210986 284294
rect 211222 284058 211306 284294
rect 211542 284058 211574 284294
rect 210954 248614 211574 284058
rect 210954 248378 210986 248614
rect 211222 248378 211306 248614
rect 211542 248378 211574 248614
rect 210954 248294 211574 248378
rect 210954 248058 210986 248294
rect 211222 248058 211306 248294
rect 211542 248058 211574 248294
rect 210954 212614 211574 248058
rect 210954 212378 210986 212614
rect 211222 212378 211306 212614
rect 211542 212378 211574 212614
rect 210954 212294 211574 212378
rect 210954 212058 210986 212294
rect 211222 212058 211306 212294
rect 211542 212058 211574 212294
rect 210954 176614 211574 212058
rect 210954 176378 210986 176614
rect 211222 176378 211306 176614
rect 211542 176378 211574 176614
rect 210954 176294 211574 176378
rect 210954 176058 210986 176294
rect 211222 176058 211306 176294
rect 211542 176058 211574 176294
rect 210954 140614 211574 176058
rect 210954 140378 210986 140614
rect 211222 140378 211306 140614
rect 211542 140378 211574 140614
rect 210954 140294 211574 140378
rect 210954 140058 210986 140294
rect 211222 140058 211306 140294
rect 211542 140058 211574 140294
rect 210954 104614 211574 140058
rect 210954 104378 210986 104614
rect 211222 104378 211306 104614
rect 211542 104378 211574 104614
rect 210954 104294 211574 104378
rect 210954 104058 210986 104294
rect 211222 104058 211306 104294
rect 211542 104058 211574 104294
rect 210954 68614 211574 104058
rect 210954 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 211574 68614
rect 210954 68294 211574 68378
rect 210954 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 211574 68294
rect 210954 32614 211574 68058
rect 210954 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 211574 32614
rect 210954 32294 211574 32378
rect 210954 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 211574 32294
rect 192954 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 193574 -6106
rect 192954 -6426 193574 -6342
rect 192954 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 193574 -6426
rect 192954 -7654 193574 -6662
rect 210954 -7066 211574 32058
rect 217794 704838 218414 705830
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 543454 218414 578898
rect 217794 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 218414 543454
rect 217794 543134 218414 543218
rect 217794 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 218414 543134
rect 217794 507454 218414 542898
rect 217794 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 218414 507454
rect 217794 507134 218414 507218
rect 217794 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 218414 507134
rect 217794 471454 218414 506898
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 217794 435454 218414 470898
rect 217794 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 218414 435454
rect 217794 435134 218414 435218
rect 217794 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 218414 435134
rect 217794 399454 218414 434898
rect 217794 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 218414 399454
rect 217794 399134 218414 399218
rect 217794 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 218414 399134
rect 217794 363454 218414 398898
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 217794 327454 218414 362898
rect 217794 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 218414 327454
rect 217794 327134 218414 327218
rect 217794 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 218414 327134
rect 217794 291454 218414 326898
rect 217794 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 218414 291454
rect 217794 291134 218414 291218
rect 217794 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 218414 291134
rect 217794 255454 218414 290898
rect 217794 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 218414 255454
rect 217794 255134 218414 255218
rect 217794 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 218414 255134
rect 217794 219454 218414 254898
rect 217794 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 218414 219454
rect 217794 219134 218414 219218
rect 217794 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 218414 219134
rect 217794 183454 218414 218898
rect 217794 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 218414 183454
rect 217794 183134 218414 183218
rect 217794 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 218414 183134
rect 217794 147454 218414 182898
rect 217794 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 218414 147454
rect 217794 147134 218414 147218
rect 217794 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 218414 147134
rect 217794 111454 218414 146898
rect 217794 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 218414 111454
rect 217794 111134 218414 111218
rect 217794 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 218414 111134
rect 217794 75454 218414 110898
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 217794 39454 218414 74898
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -1894 218414 -902
rect 221514 691174 222134 706202
rect 221514 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 222134 691174
rect 221514 690854 222134 690938
rect 221514 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 222134 690854
rect 221514 655174 222134 690618
rect 221514 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 222134 655174
rect 221514 654854 222134 654938
rect 221514 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 222134 654854
rect 221514 619174 222134 654618
rect 221514 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 222134 619174
rect 221514 618854 222134 618938
rect 221514 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 222134 618854
rect 221514 583174 222134 618618
rect 221514 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 222134 583174
rect 221514 582854 222134 582938
rect 221514 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 222134 582854
rect 221514 547174 222134 582618
rect 221514 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 222134 547174
rect 221514 546854 222134 546938
rect 221514 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 222134 546854
rect 221514 511174 222134 546618
rect 221514 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 222134 511174
rect 221514 510854 222134 510938
rect 221514 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 222134 510854
rect 221514 475174 222134 510618
rect 221514 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 222134 475174
rect 221514 474854 222134 474938
rect 221514 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 222134 474854
rect 221514 439174 222134 474618
rect 221514 438938 221546 439174
rect 221782 438938 221866 439174
rect 222102 438938 222134 439174
rect 221514 438854 222134 438938
rect 221514 438618 221546 438854
rect 221782 438618 221866 438854
rect 222102 438618 222134 438854
rect 221514 403174 222134 438618
rect 221514 402938 221546 403174
rect 221782 402938 221866 403174
rect 222102 402938 222134 403174
rect 221514 402854 222134 402938
rect 221514 402618 221546 402854
rect 221782 402618 221866 402854
rect 222102 402618 222134 402854
rect 221514 367174 222134 402618
rect 221514 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 222134 367174
rect 221514 366854 222134 366938
rect 221514 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 222134 366854
rect 221514 331174 222134 366618
rect 221514 330938 221546 331174
rect 221782 330938 221866 331174
rect 222102 330938 222134 331174
rect 221514 330854 222134 330938
rect 221514 330618 221546 330854
rect 221782 330618 221866 330854
rect 222102 330618 222134 330854
rect 221514 295174 222134 330618
rect 221514 294938 221546 295174
rect 221782 294938 221866 295174
rect 222102 294938 222134 295174
rect 221514 294854 222134 294938
rect 221514 294618 221546 294854
rect 221782 294618 221866 294854
rect 222102 294618 222134 294854
rect 221514 259174 222134 294618
rect 221514 258938 221546 259174
rect 221782 258938 221866 259174
rect 222102 258938 222134 259174
rect 221514 258854 222134 258938
rect 221514 258618 221546 258854
rect 221782 258618 221866 258854
rect 222102 258618 222134 258854
rect 221514 223174 222134 258618
rect 221514 222938 221546 223174
rect 221782 222938 221866 223174
rect 222102 222938 222134 223174
rect 221514 222854 222134 222938
rect 221514 222618 221546 222854
rect 221782 222618 221866 222854
rect 222102 222618 222134 222854
rect 221514 187174 222134 222618
rect 221514 186938 221546 187174
rect 221782 186938 221866 187174
rect 222102 186938 222134 187174
rect 221514 186854 222134 186938
rect 221514 186618 221546 186854
rect 221782 186618 221866 186854
rect 222102 186618 222134 186854
rect 221514 151174 222134 186618
rect 221514 150938 221546 151174
rect 221782 150938 221866 151174
rect 222102 150938 222134 151174
rect 221514 150854 222134 150938
rect 221514 150618 221546 150854
rect 221782 150618 221866 150854
rect 222102 150618 222134 150854
rect 221514 115174 222134 150618
rect 221514 114938 221546 115174
rect 221782 114938 221866 115174
rect 222102 114938 222134 115174
rect 221514 114854 222134 114938
rect 221514 114618 221546 114854
rect 221782 114618 221866 114854
rect 222102 114618 222134 114854
rect 221514 79174 222134 114618
rect 221514 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 222134 79174
rect 221514 78854 222134 78938
rect 221514 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 222134 78854
rect 221514 43174 222134 78618
rect 221514 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 222134 43174
rect 221514 42854 222134 42938
rect 221514 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 222134 42854
rect 221514 7174 222134 42618
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -2266 222134 6618
rect 221514 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 222134 -2266
rect 221514 -2586 222134 -2502
rect 221514 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 222134 -2586
rect 221514 -3814 222134 -2822
rect 225234 694894 225854 708122
rect 225234 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 225854 694894
rect 225234 694574 225854 694658
rect 225234 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 225854 694574
rect 225234 658894 225854 694338
rect 225234 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 225854 658894
rect 225234 658574 225854 658658
rect 225234 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 225854 658574
rect 225234 622894 225854 658338
rect 225234 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 225854 622894
rect 225234 622574 225854 622658
rect 225234 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 225854 622574
rect 225234 586894 225854 622338
rect 225234 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 225854 586894
rect 225234 586574 225854 586658
rect 225234 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 225854 586574
rect 225234 550894 225854 586338
rect 225234 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 225854 550894
rect 225234 550574 225854 550658
rect 225234 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 225854 550574
rect 225234 514894 225854 550338
rect 225234 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 225854 514894
rect 225234 514574 225854 514658
rect 225234 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 225854 514574
rect 225234 478894 225854 514338
rect 225234 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 225854 478894
rect 225234 478574 225854 478658
rect 225234 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 225854 478574
rect 225234 442894 225854 478338
rect 225234 442658 225266 442894
rect 225502 442658 225586 442894
rect 225822 442658 225854 442894
rect 225234 442574 225854 442658
rect 225234 442338 225266 442574
rect 225502 442338 225586 442574
rect 225822 442338 225854 442574
rect 225234 406894 225854 442338
rect 225234 406658 225266 406894
rect 225502 406658 225586 406894
rect 225822 406658 225854 406894
rect 225234 406574 225854 406658
rect 225234 406338 225266 406574
rect 225502 406338 225586 406574
rect 225822 406338 225854 406574
rect 225234 370894 225854 406338
rect 225234 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 225854 370894
rect 225234 370574 225854 370658
rect 225234 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 225854 370574
rect 225234 334894 225854 370338
rect 225234 334658 225266 334894
rect 225502 334658 225586 334894
rect 225822 334658 225854 334894
rect 225234 334574 225854 334658
rect 225234 334338 225266 334574
rect 225502 334338 225586 334574
rect 225822 334338 225854 334574
rect 225234 298894 225854 334338
rect 225234 298658 225266 298894
rect 225502 298658 225586 298894
rect 225822 298658 225854 298894
rect 225234 298574 225854 298658
rect 225234 298338 225266 298574
rect 225502 298338 225586 298574
rect 225822 298338 225854 298574
rect 225234 262894 225854 298338
rect 225234 262658 225266 262894
rect 225502 262658 225586 262894
rect 225822 262658 225854 262894
rect 225234 262574 225854 262658
rect 225234 262338 225266 262574
rect 225502 262338 225586 262574
rect 225822 262338 225854 262574
rect 225234 226894 225854 262338
rect 225234 226658 225266 226894
rect 225502 226658 225586 226894
rect 225822 226658 225854 226894
rect 225234 226574 225854 226658
rect 225234 226338 225266 226574
rect 225502 226338 225586 226574
rect 225822 226338 225854 226574
rect 225234 190894 225854 226338
rect 225234 190658 225266 190894
rect 225502 190658 225586 190894
rect 225822 190658 225854 190894
rect 225234 190574 225854 190658
rect 225234 190338 225266 190574
rect 225502 190338 225586 190574
rect 225822 190338 225854 190574
rect 225234 154894 225854 190338
rect 225234 154658 225266 154894
rect 225502 154658 225586 154894
rect 225822 154658 225854 154894
rect 225234 154574 225854 154658
rect 225234 154338 225266 154574
rect 225502 154338 225586 154574
rect 225822 154338 225854 154574
rect 225234 118894 225854 154338
rect 225234 118658 225266 118894
rect 225502 118658 225586 118894
rect 225822 118658 225854 118894
rect 225234 118574 225854 118658
rect 225234 118338 225266 118574
rect 225502 118338 225586 118574
rect 225822 118338 225854 118574
rect 225234 82894 225854 118338
rect 225234 82658 225266 82894
rect 225502 82658 225586 82894
rect 225822 82658 225854 82894
rect 225234 82574 225854 82658
rect 225234 82338 225266 82574
rect 225502 82338 225586 82574
rect 225822 82338 225854 82574
rect 225234 46894 225854 82338
rect 225234 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 225854 46894
rect 225234 46574 225854 46658
rect 225234 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 225854 46574
rect 225234 10894 225854 46338
rect 225234 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 225854 10894
rect 225234 10574 225854 10658
rect 225234 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 225854 10574
rect 225234 -4186 225854 10338
rect 225234 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 225854 -4186
rect 225234 -4506 225854 -4422
rect 225234 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 225854 -4506
rect 225234 -5734 225854 -4742
rect 228954 698614 229574 710042
rect 246954 711558 247574 711590
rect 246954 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 247574 711558
rect 246954 711238 247574 711322
rect 246954 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 247574 711238
rect 243234 709638 243854 709670
rect 243234 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 243854 709638
rect 243234 709318 243854 709402
rect 243234 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 243854 709318
rect 239514 707718 240134 707750
rect 239514 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 240134 707718
rect 239514 707398 240134 707482
rect 239514 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 240134 707398
rect 228954 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 229574 698614
rect 228954 698294 229574 698378
rect 228954 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 229574 698294
rect 228954 662614 229574 698058
rect 228954 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 229574 662614
rect 228954 662294 229574 662378
rect 228954 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 229574 662294
rect 228954 626614 229574 662058
rect 228954 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 229574 626614
rect 228954 626294 229574 626378
rect 228954 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 229574 626294
rect 228954 590614 229574 626058
rect 228954 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 229574 590614
rect 228954 590294 229574 590378
rect 228954 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 229574 590294
rect 228954 554614 229574 590058
rect 228954 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 229574 554614
rect 228954 554294 229574 554378
rect 228954 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 229574 554294
rect 228954 518614 229574 554058
rect 228954 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 229574 518614
rect 228954 518294 229574 518378
rect 228954 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 229574 518294
rect 228954 482614 229574 518058
rect 228954 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 229574 482614
rect 228954 482294 229574 482378
rect 228954 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 229574 482294
rect 228954 446614 229574 482058
rect 228954 446378 228986 446614
rect 229222 446378 229306 446614
rect 229542 446378 229574 446614
rect 228954 446294 229574 446378
rect 228954 446058 228986 446294
rect 229222 446058 229306 446294
rect 229542 446058 229574 446294
rect 228954 410614 229574 446058
rect 228954 410378 228986 410614
rect 229222 410378 229306 410614
rect 229542 410378 229574 410614
rect 228954 410294 229574 410378
rect 228954 410058 228986 410294
rect 229222 410058 229306 410294
rect 229542 410058 229574 410294
rect 228954 374614 229574 410058
rect 228954 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 229574 374614
rect 228954 374294 229574 374378
rect 228954 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 229574 374294
rect 228954 338614 229574 374058
rect 235794 705798 236414 705830
rect 235794 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 236414 705798
rect 235794 705478 236414 705562
rect 235794 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 236414 705478
rect 235794 669454 236414 705242
rect 239259 700364 239325 700365
rect 239259 700300 239260 700364
rect 239324 700300 239325 700364
rect 239259 700299 239325 700300
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 561454 236414 596898
rect 235794 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 236414 561454
rect 235794 561134 236414 561218
rect 235794 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 236414 561134
rect 235794 525454 236414 560898
rect 235794 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 236414 525454
rect 235794 525134 236414 525218
rect 235794 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 236414 525134
rect 235794 489454 236414 524898
rect 235794 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 236414 489454
rect 235794 489134 236414 489218
rect 235794 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 236414 489134
rect 235794 453454 236414 488898
rect 237971 466172 238037 466173
rect 237971 466108 237972 466172
rect 238036 466108 238037 466172
rect 237971 466107 238037 466108
rect 235794 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 236414 453454
rect 235794 453134 236414 453218
rect 235794 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 236414 453134
rect 235794 417454 236414 452898
rect 235794 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 236414 417454
rect 235794 417134 236414 417218
rect 235794 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 236414 417134
rect 235794 381454 236414 416898
rect 235794 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 236414 381454
rect 235794 381134 236414 381218
rect 235794 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 236414 381134
rect 235794 345454 236414 380898
rect 235794 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 236414 345454
rect 235794 345134 236414 345218
rect 235211 345132 235277 345133
rect 235211 345068 235212 345132
rect 235276 345068 235277 345132
rect 235211 345067 235277 345068
rect 228954 338378 228986 338614
rect 229222 338378 229306 338614
rect 229542 338378 229574 338614
rect 228954 338294 229574 338378
rect 228954 338058 228986 338294
rect 229222 338058 229306 338294
rect 229542 338058 229574 338294
rect 228954 302614 229574 338058
rect 228954 302378 228986 302614
rect 229222 302378 229306 302614
rect 229542 302378 229574 302614
rect 228954 302294 229574 302378
rect 228954 302058 228986 302294
rect 229222 302058 229306 302294
rect 229542 302058 229574 302294
rect 228954 266614 229574 302058
rect 228954 266378 228986 266614
rect 229222 266378 229306 266614
rect 229542 266378 229574 266614
rect 228954 266294 229574 266378
rect 228954 266058 228986 266294
rect 229222 266058 229306 266294
rect 229542 266058 229574 266294
rect 228954 230614 229574 266058
rect 228954 230378 228986 230614
rect 229222 230378 229306 230614
rect 229542 230378 229574 230614
rect 228954 230294 229574 230378
rect 228954 230058 228986 230294
rect 229222 230058 229306 230294
rect 229542 230058 229574 230294
rect 228954 194614 229574 230058
rect 228954 194378 228986 194614
rect 229222 194378 229306 194614
rect 229542 194378 229574 194614
rect 228954 194294 229574 194378
rect 228954 194058 228986 194294
rect 229222 194058 229306 194294
rect 229542 194058 229574 194294
rect 228954 158614 229574 194058
rect 235214 179349 235274 345067
rect 235794 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 236414 345134
rect 235794 309454 236414 344898
rect 237974 316029 238034 466107
rect 238523 465492 238589 465493
rect 238523 465428 238524 465492
rect 238588 465428 238589 465492
rect 238523 465427 238589 465428
rect 238339 465356 238405 465357
rect 238339 465292 238340 465356
rect 238404 465292 238405 465356
rect 238339 465291 238405 465292
rect 238155 461548 238221 461549
rect 238155 461484 238156 461548
rect 238220 461484 238221 461548
rect 238155 461483 238221 461484
rect 238158 329765 238218 461483
rect 238342 351933 238402 465291
rect 238526 356693 238586 465427
rect 238523 356692 238589 356693
rect 238523 356628 238524 356692
rect 238588 356628 238589 356692
rect 238523 356627 238589 356628
rect 238339 351932 238405 351933
rect 238339 351868 238340 351932
rect 238404 351868 238405 351932
rect 238339 351867 238405 351868
rect 238155 329764 238221 329765
rect 238155 329700 238156 329764
rect 238220 329700 238221 329764
rect 238155 329699 238221 329700
rect 237971 316028 238037 316029
rect 237971 315964 237972 316028
rect 238036 315964 238037 316028
rect 237971 315963 238037 315964
rect 235794 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 236414 309454
rect 235794 309134 236414 309218
rect 235794 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 236414 309134
rect 235579 290460 235645 290461
rect 235579 290396 235580 290460
rect 235644 290396 235645 290460
rect 235579 290395 235645 290396
rect 235395 286108 235461 286109
rect 235395 286044 235396 286108
rect 235460 286044 235461 286108
rect 235395 286043 235461 286044
rect 235398 187237 235458 286043
rect 235582 197029 235642 290395
rect 235794 273454 236414 308898
rect 235794 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 236414 273454
rect 235794 273134 236414 273218
rect 235794 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 236414 273134
rect 235794 237454 236414 272898
rect 237971 269924 238037 269925
rect 237971 269860 237972 269924
rect 238036 269860 238037 269924
rect 237971 269859 238037 269860
rect 235794 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 236414 237454
rect 235794 237134 236414 237218
rect 235794 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 236414 237134
rect 235794 201454 236414 236898
rect 235794 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 236414 201454
rect 235794 201134 236414 201218
rect 235794 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 236414 201134
rect 235579 197028 235645 197029
rect 235579 196964 235580 197028
rect 235644 196964 235645 197028
rect 235579 196963 235645 196964
rect 235395 187236 235461 187237
rect 235395 187172 235396 187236
rect 235460 187172 235461 187236
rect 235395 187171 235461 187172
rect 235211 179348 235277 179349
rect 235211 179284 235212 179348
rect 235276 179284 235277 179348
rect 235211 179283 235277 179284
rect 228954 158378 228986 158614
rect 229222 158378 229306 158614
rect 229542 158378 229574 158614
rect 228954 158294 229574 158378
rect 228954 158058 228986 158294
rect 229222 158058 229306 158294
rect 229542 158058 229574 158294
rect 228954 122614 229574 158058
rect 228954 122378 228986 122614
rect 229222 122378 229306 122614
rect 229542 122378 229574 122614
rect 228954 122294 229574 122378
rect 228954 122058 228986 122294
rect 229222 122058 229306 122294
rect 229542 122058 229574 122294
rect 228954 86614 229574 122058
rect 228954 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 229574 86614
rect 228954 86294 229574 86378
rect 228954 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 229574 86294
rect 228954 50614 229574 86058
rect 228954 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 229574 50614
rect 228954 50294 229574 50378
rect 228954 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 229574 50294
rect 228954 14614 229574 50058
rect 228954 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 229574 14614
rect 228954 14294 229574 14378
rect 228954 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 229574 14294
rect 210954 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 211574 -7066
rect 210954 -7386 211574 -7302
rect 210954 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 211574 -7386
rect 210954 -7654 211574 -7622
rect 228954 -6106 229574 14058
rect 235794 165454 236414 200898
rect 237974 199341 238034 269859
rect 238155 267340 238221 267341
rect 238155 267276 238156 267340
rect 238220 267276 238221 267340
rect 238155 267275 238221 267276
rect 237971 199340 238037 199341
rect 237971 199276 237972 199340
rect 238036 199276 238037 199340
rect 237971 199275 238037 199276
rect 238158 197573 238218 267275
rect 238339 264212 238405 264213
rect 238339 264148 238340 264212
rect 238404 264148 238405 264212
rect 238339 264147 238405 264148
rect 238155 197572 238221 197573
rect 238155 197508 238156 197572
rect 238220 197508 238221 197572
rect 238155 197507 238221 197508
rect 238342 197165 238402 264147
rect 238523 216748 238589 216749
rect 238523 216684 238524 216748
rect 238588 216684 238589 216748
rect 238523 216683 238589 216684
rect 238526 199885 238586 216683
rect 238523 199884 238589 199885
rect 238523 199820 238524 199884
rect 238588 199820 238589 199884
rect 238523 199819 238589 199820
rect 238339 197164 238405 197165
rect 238339 197100 238340 197164
rect 238404 197100 238405 197164
rect 238339 197099 238405 197100
rect 239262 179077 239322 700299
rect 239514 673174 240134 707162
rect 239514 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 240134 673174
rect 239514 672854 240134 672938
rect 239514 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 240134 672854
rect 239514 637174 240134 672618
rect 239514 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 240134 637174
rect 239514 636854 240134 636938
rect 239514 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 240134 636854
rect 239514 601174 240134 636618
rect 239514 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 240134 601174
rect 239514 600854 240134 600938
rect 239514 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 240134 600854
rect 239514 565174 240134 600618
rect 239514 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 240134 565174
rect 239514 564854 240134 564938
rect 239514 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 240134 564854
rect 239514 529174 240134 564618
rect 239514 528938 239546 529174
rect 239782 528938 239866 529174
rect 240102 528938 240134 529174
rect 239514 528854 240134 528938
rect 239514 528618 239546 528854
rect 239782 528618 239866 528854
rect 240102 528618 240134 528854
rect 239514 493174 240134 528618
rect 239514 492938 239546 493174
rect 239782 492938 239866 493174
rect 240102 492938 240134 493174
rect 239514 492854 240134 492938
rect 239514 492618 239546 492854
rect 239782 492618 239866 492854
rect 240102 492618 240134 492854
rect 239514 457174 240134 492618
rect 239514 456938 239546 457174
rect 239782 456938 239866 457174
rect 240102 456938 240134 457174
rect 239514 456854 240134 456938
rect 239514 456618 239546 456854
rect 239782 456618 239866 456854
rect 240102 456618 240134 456854
rect 239514 442000 240134 456618
rect 243234 676894 243854 709082
rect 243234 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 243854 676894
rect 243234 676574 243854 676658
rect 243234 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 243854 676574
rect 243234 640894 243854 676338
rect 243234 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 243854 640894
rect 243234 640574 243854 640658
rect 243234 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 243854 640574
rect 243234 604894 243854 640338
rect 243234 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 243854 604894
rect 243234 604574 243854 604658
rect 243234 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 243854 604574
rect 243234 568894 243854 604338
rect 243234 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 243854 568894
rect 243234 568574 243854 568658
rect 243234 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 243854 568574
rect 243234 532894 243854 568338
rect 243234 532658 243266 532894
rect 243502 532658 243586 532894
rect 243822 532658 243854 532894
rect 243234 532574 243854 532658
rect 243234 532338 243266 532574
rect 243502 532338 243586 532574
rect 243822 532338 243854 532574
rect 243234 496894 243854 532338
rect 243234 496658 243266 496894
rect 243502 496658 243586 496894
rect 243822 496658 243854 496894
rect 243234 496574 243854 496658
rect 243234 496338 243266 496574
rect 243502 496338 243586 496574
rect 243822 496338 243854 496574
rect 243234 460894 243854 496338
rect 243234 460658 243266 460894
rect 243502 460658 243586 460894
rect 243822 460658 243854 460894
rect 243234 460574 243854 460658
rect 243234 460338 243266 460574
rect 243502 460338 243586 460574
rect 243822 460338 243854 460574
rect 243234 442000 243854 460338
rect 246954 680614 247574 711002
rect 264954 710598 265574 711590
rect 264954 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 265574 710598
rect 264954 710278 265574 710362
rect 264954 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 265574 710278
rect 261234 708678 261854 709670
rect 261234 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 261854 708678
rect 261234 708358 261854 708442
rect 261234 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 261854 708358
rect 257514 706758 258134 707750
rect 257514 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 258134 706758
rect 257514 706438 258134 706522
rect 257514 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 258134 706438
rect 246954 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 247574 680614
rect 246954 680294 247574 680378
rect 246954 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 247574 680294
rect 246954 644614 247574 680058
rect 246954 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 247574 644614
rect 246954 644294 247574 644378
rect 246954 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 247574 644294
rect 246954 608614 247574 644058
rect 246954 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 247574 608614
rect 246954 608294 247574 608378
rect 246954 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 247574 608294
rect 246954 572614 247574 608058
rect 246954 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 247574 572614
rect 246954 572294 247574 572378
rect 246954 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 247574 572294
rect 246954 536614 247574 572058
rect 246954 536378 246986 536614
rect 247222 536378 247306 536614
rect 247542 536378 247574 536614
rect 246954 536294 247574 536378
rect 246954 536058 246986 536294
rect 247222 536058 247306 536294
rect 247542 536058 247574 536294
rect 246954 500614 247574 536058
rect 246954 500378 246986 500614
rect 247222 500378 247306 500614
rect 247542 500378 247574 500614
rect 246954 500294 247574 500378
rect 246954 500058 246986 500294
rect 247222 500058 247306 500294
rect 247542 500058 247574 500294
rect 246954 464614 247574 500058
rect 246954 464378 246986 464614
rect 247222 464378 247306 464614
rect 247542 464378 247574 464614
rect 246954 464294 247574 464378
rect 246954 464058 246986 464294
rect 247222 464058 247306 464294
rect 247542 464058 247574 464294
rect 246954 442000 247574 464058
rect 253794 704838 254414 705830
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 543454 254414 578898
rect 253794 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 254414 543454
rect 253794 543134 254414 543218
rect 253794 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 254414 543134
rect 253794 507454 254414 542898
rect 253794 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 254414 507454
rect 253794 507134 254414 507218
rect 253794 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 254414 507134
rect 253794 471454 254414 506898
rect 253794 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 254414 471454
rect 253794 471134 254414 471218
rect 253794 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 254414 471134
rect 253794 442000 254414 470898
rect 257514 691174 258134 706202
rect 257514 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 258134 691174
rect 257514 690854 258134 690938
rect 257514 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 258134 690854
rect 257514 655174 258134 690618
rect 257514 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 258134 655174
rect 257514 654854 258134 654938
rect 257514 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 258134 654854
rect 257514 619174 258134 654618
rect 257514 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 258134 619174
rect 257514 618854 258134 618938
rect 257514 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 258134 618854
rect 257514 583174 258134 618618
rect 257514 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 258134 583174
rect 257514 582854 258134 582938
rect 257514 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 258134 582854
rect 257514 547174 258134 582618
rect 257514 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 258134 547174
rect 257514 546854 258134 546938
rect 257514 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 258134 546854
rect 257514 511174 258134 546618
rect 257514 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 258134 511174
rect 257514 510854 258134 510938
rect 257514 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 258134 510854
rect 257514 475174 258134 510618
rect 257514 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 258134 475174
rect 257514 474854 258134 474938
rect 257514 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 258134 474854
rect 257514 442000 258134 474618
rect 261234 694894 261854 708122
rect 261234 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 261854 694894
rect 261234 694574 261854 694658
rect 261234 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 261854 694574
rect 261234 658894 261854 694338
rect 261234 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 261854 658894
rect 261234 658574 261854 658658
rect 261234 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 261854 658574
rect 261234 622894 261854 658338
rect 261234 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 261854 622894
rect 261234 622574 261854 622658
rect 261234 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 261854 622574
rect 261234 586894 261854 622338
rect 261234 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 261854 586894
rect 261234 586574 261854 586658
rect 261234 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 261854 586574
rect 261234 550894 261854 586338
rect 261234 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 261854 550894
rect 261234 550574 261854 550658
rect 261234 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 261854 550574
rect 261234 514894 261854 550338
rect 261234 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 261854 514894
rect 261234 514574 261854 514658
rect 261234 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 261854 514574
rect 261234 478894 261854 514338
rect 261234 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 261854 478894
rect 261234 478574 261854 478658
rect 261234 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 261854 478574
rect 261234 442894 261854 478338
rect 261234 442658 261266 442894
rect 261502 442658 261586 442894
rect 261822 442658 261854 442894
rect 261234 442574 261854 442658
rect 261234 442338 261266 442574
rect 261502 442338 261586 442574
rect 261822 442338 261854 442574
rect 261234 442000 261854 442338
rect 264954 698614 265574 710042
rect 282954 711558 283574 711590
rect 282954 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 283574 711558
rect 282954 711238 283574 711322
rect 282954 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 283574 711238
rect 279234 709638 279854 709670
rect 279234 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 279854 709638
rect 279234 709318 279854 709402
rect 279234 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 279854 709318
rect 275514 707718 276134 707750
rect 275514 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 276134 707718
rect 275514 707398 276134 707482
rect 275514 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 276134 707398
rect 264954 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 265574 698614
rect 264954 698294 265574 698378
rect 264954 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 265574 698294
rect 264954 662614 265574 698058
rect 264954 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 265574 662614
rect 264954 662294 265574 662378
rect 264954 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 265574 662294
rect 264954 626614 265574 662058
rect 264954 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 265574 626614
rect 264954 626294 265574 626378
rect 264954 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 265574 626294
rect 264954 590614 265574 626058
rect 264954 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 265574 590614
rect 264954 590294 265574 590378
rect 264954 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 265574 590294
rect 264954 554614 265574 590058
rect 264954 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 265574 554614
rect 264954 554294 265574 554378
rect 264954 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 265574 554294
rect 264954 518614 265574 554058
rect 264954 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 265574 518614
rect 264954 518294 265574 518378
rect 264954 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 265574 518294
rect 264954 482614 265574 518058
rect 264954 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 265574 482614
rect 264954 482294 265574 482378
rect 264954 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 265574 482294
rect 264954 446614 265574 482058
rect 264954 446378 264986 446614
rect 265222 446378 265306 446614
rect 265542 446378 265574 446614
rect 264954 446294 265574 446378
rect 264954 446058 264986 446294
rect 265222 446058 265306 446294
rect 265542 446058 265574 446294
rect 264954 442000 265574 446058
rect 271794 705798 272414 705830
rect 271794 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 272414 705798
rect 271794 705478 272414 705562
rect 271794 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 272414 705478
rect 271794 669454 272414 705242
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 561454 272414 596898
rect 271794 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 272414 561454
rect 271794 561134 272414 561218
rect 271794 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 272414 561134
rect 271794 525454 272414 560898
rect 271794 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 272414 525454
rect 271794 525134 272414 525218
rect 271794 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 272414 525134
rect 271794 489454 272414 524898
rect 271794 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 272414 489454
rect 271794 489134 272414 489218
rect 271794 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 272414 489134
rect 271794 453454 272414 488898
rect 271794 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 272414 453454
rect 271794 453134 272414 453218
rect 271794 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 272414 453134
rect 271794 442000 272414 452898
rect 275514 673174 276134 707162
rect 275514 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 276134 673174
rect 275514 672854 276134 672938
rect 275514 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 276134 672854
rect 275514 637174 276134 672618
rect 275514 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 276134 637174
rect 275514 636854 276134 636938
rect 275514 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 276134 636854
rect 275514 601174 276134 636618
rect 275514 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 276134 601174
rect 275514 600854 276134 600938
rect 275514 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 276134 600854
rect 275514 565174 276134 600618
rect 275514 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 276134 565174
rect 275514 564854 276134 564938
rect 275514 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 276134 564854
rect 275514 529174 276134 564618
rect 275514 528938 275546 529174
rect 275782 528938 275866 529174
rect 276102 528938 276134 529174
rect 275514 528854 276134 528938
rect 275514 528618 275546 528854
rect 275782 528618 275866 528854
rect 276102 528618 276134 528854
rect 275514 493174 276134 528618
rect 275514 492938 275546 493174
rect 275782 492938 275866 493174
rect 276102 492938 276134 493174
rect 275514 492854 276134 492938
rect 275514 492618 275546 492854
rect 275782 492618 275866 492854
rect 276102 492618 276134 492854
rect 275514 457174 276134 492618
rect 275514 456938 275546 457174
rect 275782 456938 275866 457174
rect 276102 456938 276134 457174
rect 275514 456854 276134 456938
rect 275514 456618 275546 456854
rect 275782 456618 275866 456854
rect 276102 456618 276134 456854
rect 275514 442000 276134 456618
rect 279234 676894 279854 709082
rect 279234 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 279854 676894
rect 279234 676574 279854 676658
rect 279234 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 279854 676574
rect 279234 640894 279854 676338
rect 279234 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 279854 640894
rect 279234 640574 279854 640658
rect 279234 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 279854 640574
rect 279234 604894 279854 640338
rect 279234 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 279854 604894
rect 279234 604574 279854 604658
rect 279234 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 279854 604574
rect 279234 568894 279854 604338
rect 279234 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 279854 568894
rect 279234 568574 279854 568658
rect 279234 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 279854 568574
rect 279234 532894 279854 568338
rect 279234 532658 279266 532894
rect 279502 532658 279586 532894
rect 279822 532658 279854 532894
rect 279234 532574 279854 532658
rect 279234 532338 279266 532574
rect 279502 532338 279586 532574
rect 279822 532338 279854 532574
rect 279234 496894 279854 532338
rect 279234 496658 279266 496894
rect 279502 496658 279586 496894
rect 279822 496658 279854 496894
rect 279234 496574 279854 496658
rect 279234 496338 279266 496574
rect 279502 496338 279586 496574
rect 279822 496338 279854 496574
rect 279234 460894 279854 496338
rect 279234 460658 279266 460894
rect 279502 460658 279586 460894
rect 279822 460658 279854 460894
rect 279234 460574 279854 460658
rect 279234 460338 279266 460574
rect 279502 460338 279586 460574
rect 279822 460338 279854 460574
rect 279234 442000 279854 460338
rect 282954 680614 283574 711002
rect 300954 710598 301574 711590
rect 300954 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 301574 710598
rect 300954 710278 301574 710362
rect 300954 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 301574 710278
rect 297234 708678 297854 709670
rect 297234 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 297854 708678
rect 297234 708358 297854 708442
rect 297234 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 297854 708358
rect 293514 706758 294134 707750
rect 293514 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 294134 706758
rect 293514 706438 294134 706522
rect 293514 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 294134 706438
rect 282954 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 283574 680614
rect 282954 680294 283574 680378
rect 282954 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 283574 680294
rect 282954 644614 283574 680058
rect 282954 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 283574 644614
rect 282954 644294 283574 644378
rect 282954 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 283574 644294
rect 282954 608614 283574 644058
rect 282954 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 283574 608614
rect 282954 608294 283574 608378
rect 282954 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 283574 608294
rect 282954 572614 283574 608058
rect 282954 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 283574 572614
rect 282954 572294 283574 572378
rect 282954 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 283574 572294
rect 282954 536614 283574 572058
rect 282954 536378 282986 536614
rect 283222 536378 283306 536614
rect 283542 536378 283574 536614
rect 282954 536294 283574 536378
rect 282954 536058 282986 536294
rect 283222 536058 283306 536294
rect 283542 536058 283574 536294
rect 282954 500614 283574 536058
rect 282954 500378 282986 500614
rect 283222 500378 283306 500614
rect 283542 500378 283574 500614
rect 282954 500294 283574 500378
rect 282954 500058 282986 500294
rect 283222 500058 283306 500294
rect 283542 500058 283574 500294
rect 282954 464614 283574 500058
rect 282954 464378 282986 464614
rect 283222 464378 283306 464614
rect 283542 464378 283574 464614
rect 282954 464294 283574 464378
rect 282954 464058 282986 464294
rect 283222 464058 283306 464294
rect 283542 464058 283574 464294
rect 282954 442000 283574 464058
rect 289794 704838 290414 705830
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 543454 290414 578898
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289794 507454 290414 542898
rect 289794 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 290414 507454
rect 289794 507134 290414 507218
rect 289794 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 290414 507134
rect 289794 471454 290414 506898
rect 289794 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 290414 471454
rect 289794 471134 290414 471218
rect 289794 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 290414 471134
rect 289794 442000 290414 470898
rect 293514 691174 294134 706202
rect 293514 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 294134 691174
rect 293514 690854 294134 690938
rect 293514 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 294134 690854
rect 293514 655174 294134 690618
rect 293514 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 294134 655174
rect 293514 654854 294134 654938
rect 293514 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 294134 654854
rect 293514 619174 294134 654618
rect 293514 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 294134 619174
rect 293514 618854 294134 618938
rect 293514 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 294134 618854
rect 293514 583174 294134 618618
rect 293514 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 294134 583174
rect 293514 582854 294134 582938
rect 293514 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 294134 582854
rect 293514 547174 294134 582618
rect 293514 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 294134 547174
rect 293514 546854 294134 546938
rect 293514 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 294134 546854
rect 293514 511174 294134 546618
rect 293514 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 294134 511174
rect 293514 510854 294134 510938
rect 293514 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 294134 510854
rect 293514 475174 294134 510618
rect 293514 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 294134 475174
rect 293514 474854 294134 474938
rect 293514 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 294134 474854
rect 293514 442000 294134 474618
rect 297234 694894 297854 708122
rect 297234 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 297854 694894
rect 297234 694574 297854 694658
rect 297234 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 297854 694574
rect 297234 658894 297854 694338
rect 297234 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 297854 658894
rect 297234 658574 297854 658658
rect 297234 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 297854 658574
rect 297234 622894 297854 658338
rect 297234 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 297854 622894
rect 297234 622574 297854 622658
rect 297234 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 297854 622574
rect 297234 586894 297854 622338
rect 297234 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 297854 586894
rect 297234 586574 297854 586658
rect 297234 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 297854 586574
rect 297234 550894 297854 586338
rect 297234 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 297854 550894
rect 297234 550574 297854 550658
rect 297234 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 297854 550574
rect 297234 514894 297854 550338
rect 297234 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 297854 514894
rect 297234 514574 297854 514658
rect 297234 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 297854 514574
rect 297234 478894 297854 514338
rect 297234 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 297854 478894
rect 297234 478574 297854 478658
rect 297234 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 297854 478574
rect 297234 442894 297854 478338
rect 297234 442658 297266 442894
rect 297502 442658 297586 442894
rect 297822 442658 297854 442894
rect 297234 442574 297854 442658
rect 297234 442338 297266 442574
rect 297502 442338 297586 442574
rect 297822 442338 297854 442574
rect 297234 442000 297854 442338
rect 300954 698614 301574 710042
rect 318954 711558 319574 711590
rect 318954 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 319574 711558
rect 318954 711238 319574 711322
rect 318954 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 319574 711238
rect 315234 709638 315854 709670
rect 315234 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 315854 709638
rect 315234 709318 315854 709402
rect 315234 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 315854 709318
rect 311514 707718 312134 707750
rect 311514 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 312134 707718
rect 311514 707398 312134 707482
rect 311514 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 312134 707398
rect 300954 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 301574 698614
rect 300954 698294 301574 698378
rect 300954 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 301574 698294
rect 300954 662614 301574 698058
rect 300954 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 301574 662614
rect 300954 662294 301574 662378
rect 300954 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 301574 662294
rect 300954 626614 301574 662058
rect 300954 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 301574 626614
rect 300954 626294 301574 626378
rect 300954 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 301574 626294
rect 300954 590614 301574 626058
rect 300954 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 301574 590614
rect 300954 590294 301574 590378
rect 300954 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 301574 590294
rect 300954 554614 301574 590058
rect 300954 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 301574 554614
rect 300954 554294 301574 554378
rect 300954 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 301574 554294
rect 300954 518614 301574 554058
rect 300954 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 301574 518614
rect 300954 518294 301574 518378
rect 300954 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 301574 518294
rect 300954 482614 301574 518058
rect 300954 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 301574 482614
rect 300954 482294 301574 482378
rect 300954 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 301574 482294
rect 300954 446614 301574 482058
rect 300954 446378 300986 446614
rect 301222 446378 301306 446614
rect 301542 446378 301574 446614
rect 300954 446294 301574 446378
rect 300954 446058 300986 446294
rect 301222 446058 301306 446294
rect 301542 446058 301574 446294
rect 300954 442000 301574 446058
rect 307794 705798 308414 705830
rect 307794 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 308414 705798
rect 307794 705478 308414 705562
rect 307794 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 308414 705478
rect 307794 669454 308414 705242
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 561454 308414 596898
rect 307794 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 308414 561454
rect 307794 561134 308414 561218
rect 307794 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 308414 561134
rect 307794 525454 308414 560898
rect 307794 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 308414 525454
rect 307794 525134 308414 525218
rect 307794 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 308414 525134
rect 307794 489454 308414 524898
rect 307794 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 308414 489454
rect 307794 489134 308414 489218
rect 307794 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 308414 489134
rect 307794 453454 308414 488898
rect 307794 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 308414 453454
rect 307794 453134 308414 453218
rect 307794 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 308414 453134
rect 307794 442000 308414 452898
rect 311514 673174 312134 707162
rect 311514 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 312134 673174
rect 311514 672854 312134 672938
rect 311514 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 312134 672854
rect 311514 637174 312134 672618
rect 311514 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 312134 637174
rect 311514 636854 312134 636938
rect 311514 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 312134 636854
rect 311514 601174 312134 636618
rect 311514 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 312134 601174
rect 311514 600854 312134 600938
rect 311514 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 312134 600854
rect 311514 565174 312134 600618
rect 311514 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 312134 565174
rect 311514 564854 312134 564938
rect 311514 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 312134 564854
rect 311514 529174 312134 564618
rect 311514 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 312134 529174
rect 311514 528854 312134 528938
rect 311514 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 312134 528854
rect 311514 493174 312134 528618
rect 311514 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 312134 493174
rect 311514 492854 312134 492938
rect 311514 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 312134 492854
rect 311514 457174 312134 492618
rect 311514 456938 311546 457174
rect 311782 456938 311866 457174
rect 312102 456938 312134 457174
rect 311514 456854 312134 456938
rect 311514 456618 311546 456854
rect 311782 456618 311866 456854
rect 312102 456618 312134 456854
rect 311514 442000 312134 456618
rect 315234 676894 315854 709082
rect 315234 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 315854 676894
rect 315234 676574 315854 676658
rect 315234 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 315854 676574
rect 315234 640894 315854 676338
rect 315234 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 315854 640894
rect 315234 640574 315854 640658
rect 315234 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 315854 640574
rect 315234 604894 315854 640338
rect 315234 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 315854 604894
rect 315234 604574 315854 604658
rect 315234 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 315854 604574
rect 315234 568894 315854 604338
rect 315234 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 315854 568894
rect 315234 568574 315854 568658
rect 315234 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 315854 568574
rect 315234 532894 315854 568338
rect 315234 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 315854 532894
rect 315234 532574 315854 532658
rect 315234 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 315854 532574
rect 315234 496894 315854 532338
rect 315234 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 315854 496894
rect 315234 496574 315854 496658
rect 315234 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 315854 496574
rect 315234 460894 315854 496338
rect 315234 460658 315266 460894
rect 315502 460658 315586 460894
rect 315822 460658 315854 460894
rect 315234 460574 315854 460658
rect 315234 460338 315266 460574
rect 315502 460338 315586 460574
rect 315822 460338 315854 460574
rect 315234 442000 315854 460338
rect 318954 680614 319574 711002
rect 336954 710598 337574 711590
rect 336954 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 337574 710598
rect 336954 710278 337574 710362
rect 336954 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 337574 710278
rect 333234 708678 333854 709670
rect 333234 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 333854 708678
rect 333234 708358 333854 708442
rect 333234 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 333854 708358
rect 329514 706758 330134 707750
rect 329514 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 330134 706758
rect 329514 706438 330134 706522
rect 329514 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 330134 706438
rect 318954 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 319574 680614
rect 318954 680294 319574 680378
rect 318954 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 319574 680294
rect 318954 644614 319574 680058
rect 318954 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 319574 644614
rect 318954 644294 319574 644378
rect 318954 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 319574 644294
rect 318954 608614 319574 644058
rect 318954 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 319574 608614
rect 318954 608294 319574 608378
rect 318954 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 319574 608294
rect 318954 572614 319574 608058
rect 318954 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 319574 572614
rect 318954 572294 319574 572378
rect 318954 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 319574 572294
rect 318954 536614 319574 572058
rect 318954 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 319574 536614
rect 318954 536294 319574 536378
rect 318954 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 319574 536294
rect 318954 500614 319574 536058
rect 318954 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 319574 500614
rect 318954 500294 319574 500378
rect 318954 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 319574 500294
rect 318954 464614 319574 500058
rect 318954 464378 318986 464614
rect 319222 464378 319306 464614
rect 319542 464378 319574 464614
rect 318954 464294 319574 464378
rect 318954 464058 318986 464294
rect 319222 464058 319306 464294
rect 319542 464058 319574 464294
rect 318954 442000 319574 464058
rect 325794 704838 326414 705830
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 543454 326414 578898
rect 325794 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 326414 543454
rect 325794 543134 326414 543218
rect 325794 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 326414 543134
rect 325794 507454 326414 542898
rect 325794 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 326414 507454
rect 325794 507134 326414 507218
rect 325794 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 326414 507134
rect 325794 471454 326414 506898
rect 325794 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 326414 471454
rect 325794 471134 326414 471218
rect 325794 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 326414 471134
rect 325794 442000 326414 470898
rect 329514 691174 330134 706202
rect 329514 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 330134 691174
rect 329514 690854 330134 690938
rect 329514 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 330134 690854
rect 329514 655174 330134 690618
rect 329514 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 330134 655174
rect 329514 654854 330134 654938
rect 329514 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 330134 654854
rect 329514 619174 330134 654618
rect 329514 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 330134 619174
rect 329514 618854 330134 618938
rect 329514 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 330134 618854
rect 329514 583174 330134 618618
rect 329514 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 330134 583174
rect 329514 582854 330134 582938
rect 329514 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 330134 582854
rect 329514 547174 330134 582618
rect 329514 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 330134 547174
rect 329514 546854 330134 546938
rect 329514 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 330134 546854
rect 329514 511174 330134 546618
rect 329514 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 330134 511174
rect 329514 510854 330134 510938
rect 329514 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 330134 510854
rect 329514 475174 330134 510618
rect 329514 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 330134 475174
rect 329514 474854 330134 474938
rect 329514 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 330134 474854
rect 329514 442000 330134 474618
rect 333234 694894 333854 708122
rect 333234 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 333854 694894
rect 333234 694574 333854 694658
rect 333234 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 333854 694574
rect 333234 658894 333854 694338
rect 333234 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 333854 658894
rect 333234 658574 333854 658658
rect 333234 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 333854 658574
rect 333234 622894 333854 658338
rect 333234 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 333854 622894
rect 333234 622574 333854 622658
rect 333234 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 333854 622574
rect 333234 586894 333854 622338
rect 333234 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 333854 586894
rect 333234 586574 333854 586658
rect 333234 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 333854 586574
rect 333234 550894 333854 586338
rect 333234 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 333854 550894
rect 333234 550574 333854 550658
rect 333234 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 333854 550574
rect 333234 514894 333854 550338
rect 333234 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 333854 514894
rect 333234 514574 333854 514658
rect 333234 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 333854 514574
rect 333234 478894 333854 514338
rect 333234 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 333854 478894
rect 333234 478574 333854 478658
rect 333234 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 333854 478574
rect 333234 442894 333854 478338
rect 333234 442658 333266 442894
rect 333502 442658 333586 442894
rect 333822 442658 333854 442894
rect 333234 442574 333854 442658
rect 333234 442338 333266 442574
rect 333502 442338 333586 442574
rect 333822 442338 333854 442574
rect 333234 442000 333854 442338
rect 336954 698614 337574 710042
rect 354954 711558 355574 711590
rect 354954 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 355574 711558
rect 354954 711238 355574 711322
rect 354954 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 355574 711238
rect 351234 709638 351854 709670
rect 351234 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 351854 709638
rect 351234 709318 351854 709402
rect 351234 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 351854 709318
rect 347514 707718 348134 707750
rect 347514 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 348134 707718
rect 347514 707398 348134 707482
rect 347514 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 348134 707398
rect 336954 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 337574 698614
rect 336954 698294 337574 698378
rect 336954 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 337574 698294
rect 336954 662614 337574 698058
rect 336954 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 337574 662614
rect 336954 662294 337574 662378
rect 336954 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 337574 662294
rect 336954 626614 337574 662058
rect 336954 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 337574 626614
rect 336954 626294 337574 626378
rect 336954 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 337574 626294
rect 336954 590614 337574 626058
rect 336954 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 337574 590614
rect 336954 590294 337574 590378
rect 336954 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 337574 590294
rect 336954 554614 337574 590058
rect 336954 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 337574 554614
rect 336954 554294 337574 554378
rect 336954 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 337574 554294
rect 336954 518614 337574 554058
rect 336954 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 337574 518614
rect 336954 518294 337574 518378
rect 336954 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 337574 518294
rect 336954 482614 337574 518058
rect 336954 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 337574 482614
rect 336954 482294 337574 482378
rect 336954 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 337574 482294
rect 336954 446614 337574 482058
rect 336954 446378 336986 446614
rect 337222 446378 337306 446614
rect 337542 446378 337574 446614
rect 336954 446294 337574 446378
rect 336954 446058 336986 446294
rect 337222 446058 337306 446294
rect 337542 446058 337574 446294
rect 336954 442000 337574 446058
rect 343794 705798 344414 705830
rect 343794 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 344414 705798
rect 343794 705478 344414 705562
rect 343794 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 344414 705478
rect 343794 669454 344414 705242
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 561454 344414 596898
rect 343794 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 344414 561454
rect 343794 561134 344414 561218
rect 343794 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 344414 561134
rect 343794 525454 344414 560898
rect 343794 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 344414 525454
rect 343794 525134 344414 525218
rect 343794 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 344414 525134
rect 343794 489454 344414 524898
rect 343794 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 344414 489454
rect 343794 489134 344414 489218
rect 343794 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 344414 489134
rect 343794 453454 344414 488898
rect 343794 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 344414 453454
rect 343794 453134 344414 453218
rect 343794 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 344414 453134
rect 343794 442000 344414 452898
rect 347514 673174 348134 707162
rect 347514 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 348134 673174
rect 347514 672854 348134 672938
rect 347514 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 348134 672854
rect 347514 637174 348134 672618
rect 347514 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 348134 637174
rect 347514 636854 348134 636938
rect 347514 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 348134 636854
rect 347514 601174 348134 636618
rect 347514 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 348134 601174
rect 347514 600854 348134 600938
rect 347514 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 348134 600854
rect 347514 565174 348134 600618
rect 347514 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 348134 565174
rect 347514 564854 348134 564938
rect 347514 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 348134 564854
rect 347514 529174 348134 564618
rect 347514 528938 347546 529174
rect 347782 528938 347866 529174
rect 348102 528938 348134 529174
rect 347514 528854 348134 528938
rect 347514 528618 347546 528854
rect 347782 528618 347866 528854
rect 348102 528618 348134 528854
rect 347514 493174 348134 528618
rect 347514 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 348134 493174
rect 347514 492854 348134 492938
rect 347514 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 348134 492854
rect 347514 457174 348134 492618
rect 347514 456938 347546 457174
rect 347782 456938 347866 457174
rect 348102 456938 348134 457174
rect 347514 456854 348134 456938
rect 347514 456618 347546 456854
rect 347782 456618 347866 456854
rect 348102 456618 348134 456854
rect 347514 442000 348134 456618
rect 351234 676894 351854 709082
rect 351234 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 351854 676894
rect 351234 676574 351854 676658
rect 351234 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 351854 676574
rect 351234 640894 351854 676338
rect 351234 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 351854 640894
rect 351234 640574 351854 640658
rect 351234 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 351854 640574
rect 351234 604894 351854 640338
rect 351234 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 351854 604894
rect 351234 604574 351854 604658
rect 351234 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 351854 604574
rect 351234 568894 351854 604338
rect 351234 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 351854 568894
rect 351234 568574 351854 568658
rect 351234 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 351854 568574
rect 351234 532894 351854 568338
rect 351234 532658 351266 532894
rect 351502 532658 351586 532894
rect 351822 532658 351854 532894
rect 351234 532574 351854 532658
rect 351234 532338 351266 532574
rect 351502 532338 351586 532574
rect 351822 532338 351854 532574
rect 351234 496894 351854 532338
rect 351234 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 351854 496894
rect 351234 496574 351854 496658
rect 351234 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 351854 496574
rect 351234 460894 351854 496338
rect 351234 460658 351266 460894
rect 351502 460658 351586 460894
rect 351822 460658 351854 460894
rect 351234 460574 351854 460658
rect 351234 460338 351266 460574
rect 351502 460338 351586 460574
rect 351822 460338 351854 460574
rect 351234 442000 351854 460338
rect 354954 680614 355574 711002
rect 372954 710598 373574 711590
rect 372954 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 373574 710598
rect 372954 710278 373574 710362
rect 372954 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 373574 710278
rect 369234 708678 369854 709670
rect 369234 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 369854 708678
rect 369234 708358 369854 708442
rect 369234 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 369854 708358
rect 365514 706758 366134 707750
rect 365514 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 366134 706758
rect 365514 706438 366134 706522
rect 365514 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 366134 706438
rect 354954 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 355574 680614
rect 354954 680294 355574 680378
rect 354954 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 355574 680294
rect 354954 644614 355574 680058
rect 354954 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 355574 644614
rect 354954 644294 355574 644378
rect 354954 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 355574 644294
rect 354954 608614 355574 644058
rect 354954 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 355574 608614
rect 354954 608294 355574 608378
rect 354954 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 355574 608294
rect 354954 572614 355574 608058
rect 354954 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 355574 572614
rect 354954 572294 355574 572378
rect 354954 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 355574 572294
rect 354954 536614 355574 572058
rect 354954 536378 354986 536614
rect 355222 536378 355306 536614
rect 355542 536378 355574 536614
rect 354954 536294 355574 536378
rect 354954 536058 354986 536294
rect 355222 536058 355306 536294
rect 355542 536058 355574 536294
rect 354954 500614 355574 536058
rect 354954 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 355574 500614
rect 354954 500294 355574 500378
rect 354954 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 355574 500294
rect 354954 464614 355574 500058
rect 354954 464378 354986 464614
rect 355222 464378 355306 464614
rect 355542 464378 355574 464614
rect 354954 464294 355574 464378
rect 354954 464058 354986 464294
rect 355222 464058 355306 464294
rect 355542 464058 355574 464294
rect 354954 442000 355574 464058
rect 361794 704838 362414 705830
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 442000 362414 470898
rect 365514 691174 366134 706202
rect 365514 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 366134 691174
rect 365514 690854 366134 690938
rect 365514 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 366134 690854
rect 365514 655174 366134 690618
rect 365514 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 366134 655174
rect 365514 654854 366134 654938
rect 365514 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 366134 654854
rect 365514 619174 366134 654618
rect 365514 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 366134 619174
rect 365514 618854 366134 618938
rect 365514 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 366134 618854
rect 365514 583174 366134 618618
rect 365514 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 366134 583174
rect 365514 582854 366134 582938
rect 365514 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 366134 582854
rect 365514 547174 366134 582618
rect 365514 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 366134 547174
rect 365514 546854 366134 546938
rect 365514 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 366134 546854
rect 365514 511174 366134 546618
rect 365514 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 366134 511174
rect 365514 510854 366134 510938
rect 365514 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 366134 510854
rect 365514 475174 366134 510618
rect 365514 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 366134 475174
rect 365514 474854 366134 474938
rect 365514 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 366134 474854
rect 365514 442000 366134 474618
rect 369234 694894 369854 708122
rect 369234 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 369854 694894
rect 369234 694574 369854 694658
rect 369234 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 369854 694574
rect 369234 658894 369854 694338
rect 369234 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 369854 658894
rect 369234 658574 369854 658658
rect 369234 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 369854 658574
rect 369234 622894 369854 658338
rect 369234 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 369854 622894
rect 369234 622574 369854 622658
rect 369234 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 369854 622574
rect 369234 586894 369854 622338
rect 369234 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 369854 586894
rect 369234 586574 369854 586658
rect 369234 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 369854 586574
rect 369234 550894 369854 586338
rect 369234 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 369854 550894
rect 369234 550574 369854 550658
rect 369234 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 369854 550574
rect 369234 514894 369854 550338
rect 369234 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 369854 514894
rect 369234 514574 369854 514658
rect 369234 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 369854 514574
rect 369234 478894 369854 514338
rect 369234 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 369854 478894
rect 369234 478574 369854 478658
rect 369234 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 369854 478574
rect 369234 442894 369854 478338
rect 369234 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 369854 442894
rect 369234 442574 369854 442658
rect 369234 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 369854 442574
rect 369234 442000 369854 442338
rect 372954 698614 373574 710042
rect 390954 711558 391574 711590
rect 390954 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 391574 711558
rect 390954 711238 391574 711322
rect 390954 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 391574 711238
rect 387234 709638 387854 709670
rect 387234 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 387854 709638
rect 387234 709318 387854 709402
rect 387234 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 387854 709318
rect 383514 707718 384134 707750
rect 383514 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 384134 707718
rect 383514 707398 384134 707482
rect 383514 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 384134 707398
rect 372954 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 373574 698614
rect 372954 698294 373574 698378
rect 372954 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 373574 698294
rect 372954 662614 373574 698058
rect 372954 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 373574 662614
rect 372954 662294 373574 662378
rect 372954 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 373574 662294
rect 372954 626614 373574 662058
rect 372954 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 373574 626614
rect 372954 626294 373574 626378
rect 372954 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 373574 626294
rect 372954 590614 373574 626058
rect 372954 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 373574 590614
rect 372954 590294 373574 590378
rect 372954 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 373574 590294
rect 372954 554614 373574 590058
rect 372954 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 373574 554614
rect 372954 554294 373574 554378
rect 372954 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 373574 554294
rect 372954 518614 373574 554058
rect 372954 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 373574 518614
rect 372954 518294 373574 518378
rect 372954 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 373574 518294
rect 372954 482614 373574 518058
rect 372954 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 373574 482614
rect 372954 482294 373574 482378
rect 372954 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 373574 482294
rect 372954 446614 373574 482058
rect 372954 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 373574 446614
rect 372954 446294 373574 446378
rect 372954 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 373574 446294
rect 372954 442000 373574 446058
rect 379794 705798 380414 705830
rect 379794 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 380414 705798
rect 379794 705478 380414 705562
rect 379794 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 380414 705478
rect 379794 669454 380414 705242
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 561454 380414 596898
rect 379794 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 380414 561454
rect 379794 561134 380414 561218
rect 379794 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 380414 561134
rect 379794 525454 380414 560898
rect 379794 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 380414 525454
rect 379794 525134 380414 525218
rect 379794 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 380414 525134
rect 379794 489454 380414 524898
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 379794 453454 380414 488898
rect 379794 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 380414 453454
rect 379794 453134 380414 453218
rect 379794 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 380414 453134
rect 379794 442000 380414 452898
rect 383514 673174 384134 707162
rect 383514 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 384134 673174
rect 383514 672854 384134 672938
rect 383514 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 384134 672854
rect 383514 637174 384134 672618
rect 383514 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 384134 637174
rect 383514 636854 384134 636938
rect 383514 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 384134 636854
rect 383514 601174 384134 636618
rect 383514 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 384134 601174
rect 383514 600854 384134 600938
rect 383514 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 384134 600854
rect 383514 565174 384134 600618
rect 383514 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 384134 565174
rect 383514 564854 384134 564938
rect 383514 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 384134 564854
rect 383514 529174 384134 564618
rect 383514 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 384134 529174
rect 383514 528854 384134 528938
rect 383514 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 384134 528854
rect 383514 493174 384134 528618
rect 383514 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 384134 493174
rect 383514 492854 384134 492938
rect 383514 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 384134 492854
rect 383514 457174 384134 492618
rect 383514 456938 383546 457174
rect 383782 456938 383866 457174
rect 384102 456938 384134 457174
rect 383514 456854 384134 456938
rect 383514 456618 383546 456854
rect 383782 456618 383866 456854
rect 384102 456618 384134 456854
rect 383514 442000 384134 456618
rect 387234 676894 387854 709082
rect 387234 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 387854 676894
rect 387234 676574 387854 676658
rect 387234 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 387854 676574
rect 387234 640894 387854 676338
rect 387234 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 387854 640894
rect 387234 640574 387854 640658
rect 387234 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 387854 640574
rect 387234 604894 387854 640338
rect 387234 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 387854 604894
rect 387234 604574 387854 604658
rect 387234 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 387854 604574
rect 387234 568894 387854 604338
rect 387234 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 387854 568894
rect 387234 568574 387854 568658
rect 387234 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 387854 568574
rect 387234 532894 387854 568338
rect 387234 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 387854 532894
rect 387234 532574 387854 532658
rect 387234 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 387854 532574
rect 387234 496894 387854 532338
rect 387234 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 387854 496894
rect 387234 496574 387854 496658
rect 387234 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 387854 496574
rect 387234 460894 387854 496338
rect 387234 460658 387266 460894
rect 387502 460658 387586 460894
rect 387822 460658 387854 460894
rect 387234 460574 387854 460658
rect 387234 460338 387266 460574
rect 387502 460338 387586 460574
rect 387822 460338 387854 460574
rect 387234 442000 387854 460338
rect 390954 680614 391574 711002
rect 408954 710598 409574 711590
rect 408954 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 409574 710598
rect 408954 710278 409574 710362
rect 408954 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 409574 710278
rect 405234 708678 405854 709670
rect 405234 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 405854 708678
rect 405234 708358 405854 708442
rect 405234 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 405854 708358
rect 401514 706758 402134 707750
rect 401514 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 402134 706758
rect 401514 706438 402134 706522
rect 401514 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 402134 706438
rect 390954 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 391574 680614
rect 390954 680294 391574 680378
rect 390954 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 391574 680294
rect 390954 644614 391574 680058
rect 390954 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 391574 644614
rect 390954 644294 391574 644378
rect 390954 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 391574 644294
rect 390954 608614 391574 644058
rect 390954 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 391574 608614
rect 390954 608294 391574 608378
rect 390954 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 391574 608294
rect 390954 572614 391574 608058
rect 390954 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 391574 572614
rect 390954 572294 391574 572378
rect 390954 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 391574 572294
rect 390954 536614 391574 572058
rect 390954 536378 390986 536614
rect 391222 536378 391306 536614
rect 391542 536378 391574 536614
rect 390954 536294 391574 536378
rect 390954 536058 390986 536294
rect 391222 536058 391306 536294
rect 391542 536058 391574 536294
rect 390954 500614 391574 536058
rect 390954 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 391574 500614
rect 390954 500294 391574 500378
rect 390954 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 391574 500294
rect 390954 464614 391574 500058
rect 390954 464378 390986 464614
rect 391222 464378 391306 464614
rect 391542 464378 391574 464614
rect 390954 464294 391574 464378
rect 390954 464058 390986 464294
rect 391222 464058 391306 464294
rect 391542 464058 391574 464294
rect 390954 442000 391574 464058
rect 397794 704838 398414 705830
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 442000 398414 470898
rect 401514 691174 402134 706202
rect 401514 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 402134 691174
rect 401514 690854 402134 690938
rect 401514 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 402134 690854
rect 401514 655174 402134 690618
rect 401514 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 402134 655174
rect 401514 654854 402134 654938
rect 401514 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 402134 654854
rect 401514 619174 402134 654618
rect 401514 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 402134 619174
rect 401514 618854 402134 618938
rect 401514 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 402134 618854
rect 401514 583174 402134 618618
rect 401514 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 402134 583174
rect 401514 582854 402134 582938
rect 401514 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 402134 582854
rect 401514 547174 402134 582618
rect 401514 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 402134 547174
rect 401514 546854 402134 546938
rect 401514 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 402134 546854
rect 401514 511174 402134 546618
rect 401514 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 402134 511174
rect 401514 510854 402134 510938
rect 401514 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 402134 510854
rect 401514 475174 402134 510618
rect 401514 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 402134 475174
rect 401514 474854 402134 474938
rect 401514 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 402134 474854
rect 401514 442000 402134 474618
rect 405234 694894 405854 708122
rect 405234 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 405854 694894
rect 405234 694574 405854 694658
rect 405234 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 405854 694574
rect 405234 658894 405854 694338
rect 405234 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 405854 658894
rect 405234 658574 405854 658658
rect 405234 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 405854 658574
rect 405234 622894 405854 658338
rect 405234 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 405854 622894
rect 405234 622574 405854 622658
rect 405234 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 405854 622574
rect 405234 586894 405854 622338
rect 405234 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 405854 586894
rect 405234 586574 405854 586658
rect 405234 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 405854 586574
rect 405234 550894 405854 586338
rect 405234 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 405854 550894
rect 405234 550574 405854 550658
rect 405234 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 405854 550574
rect 405234 514894 405854 550338
rect 405234 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 405854 514894
rect 405234 514574 405854 514658
rect 405234 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 405854 514574
rect 405234 478894 405854 514338
rect 405234 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 405854 478894
rect 405234 478574 405854 478658
rect 405234 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 405854 478574
rect 405234 442894 405854 478338
rect 405234 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 405854 442894
rect 405234 442574 405854 442658
rect 405234 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 405854 442574
rect 405234 442000 405854 442338
rect 408954 698614 409574 710042
rect 426954 711558 427574 711590
rect 426954 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 427574 711558
rect 426954 711238 427574 711322
rect 426954 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 427574 711238
rect 423234 709638 423854 709670
rect 423234 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 423854 709638
rect 423234 709318 423854 709402
rect 423234 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 423854 709318
rect 419514 707718 420134 707750
rect 419514 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 420134 707718
rect 419514 707398 420134 707482
rect 419514 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 420134 707398
rect 408954 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 409574 698614
rect 408954 698294 409574 698378
rect 408954 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 409574 698294
rect 408954 662614 409574 698058
rect 408954 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 409574 662614
rect 408954 662294 409574 662378
rect 408954 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 409574 662294
rect 408954 626614 409574 662058
rect 408954 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 409574 626614
rect 408954 626294 409574 626378
rect 408954 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 409574 626294
rect 408954 590614 409574 626058
rect 408954 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 409574 590614
rect 408954 590294 409574 590378
rect 408954 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 409574 590294
rect 408954 554614 409574 590058
rect 408954 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 409574 554614
rect 408954 554294 409574 554378
rect 408954 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 409574 554294
rect 408954 518614 409574 554058
rect 408954 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 409574 518614
rect 408954 518294 409574 518378
rect 408954 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 409574 518294
rect 408954 482614 409574 518058
rect 408954 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 409574 482614
rect 408954 482294 409574 482378
rect 408954 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 409574 482294
rect 408954 446614 409574 482058
rect 408954 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 409574 446614
rect 408954 446294 409574 446378
rect 408954 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 409574 446294
rect 408954 442000 409574 446058
rect 415794 705798 416414 705830
rect 415794 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 416414 705798
rect 415794 705478 416414 705562
rect 415794 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 416414 705478
rect 415794 669454 416414 705242
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 561454 416414 596898
rect 415794 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 416414 561454
rect 415794 561134 416414 561218
rect 415794 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 416414 561134
rect 415794 525454 416414 560898
rect 415794 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 416414 525454
rect 415794 525134 416414 525218
rect 415794 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 416414 525134
rect 415794 489454 416414 524898
rect 415794 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 416414 489454
rect 415794 489134 416414 489218
rect 415794 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 416414 489134
rect 415794 453454 416414 488898
rect 415794 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 416414 453454
rect 415794 453134 416414 453218
rect 415794 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 416414 453134
rect 415794 442000 416414 452898
rect 419514 673174 420134 707162
rect 419514 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 420134 673174
rect 419514 672854 420134 672938
rect 419514 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 420134 672854
rect 419514 637174 420134 672618
rect 419514 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 420134 637174
rect 419514 636854 420134 636938
rect 419514 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 420134 636854
rect 419514 601174 420134 636618
rect 419514 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 420134 601174
rect 419514 600854 420134 600938
rect 419514 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 420134 600854
rect 419514 565174 420134 600618
rect 419514 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 420134 565174
rect 419514 564854 420134 564938
rect 419514 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 420134 564854
rect 419514 529174 420134 564618
rect 419514 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 420134 529174
rect 419514 528854 420134 528938
rect 419514 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 420134 528854
rect 419514 493174 420134 528618
rect 419514 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 420134 493174
rect 419514 492854 420134 492938
rect 419514 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 420134 492854
rect 419514 457174 420134 492618
rect 419514 456938 419546 457174
rect 419782 456938 419866 457174
rect 420102 456938 420134 457174
rect 419514 456854 420134 456938
rect 419514 456618 419546 456854
rect 419782 456618 419866 456854
rect 420102 456618 420134 456854
rect 419514 442000 420134 456618
rect 423234 676894 423854 709082
rect 423234 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 423854 676894
rect 423234 676574 423854 676658
rect 423234 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 423854 676574
rect 423234 640894 423854 676338
rect 423234 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 423854 640894
rect 423234 640574 423854 640658
rect 423234 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 423854 640574
rect 423234 604894 423854 640338
rect 423234 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 423854 604894
rect 423234 604574 423854 604658
rect 423234 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 423854 604574
rect 423234 568894 423854 604338
rect 423234 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 423854 568894
rect 423234 568574 423854 568658
rect 423234 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 423854 568574
rect 423234 532894 423854 568338
rect 423234 532658 423266 532894
rect 423502 532658 423586 532894
rect 423822 532658 423854 532894
rect 423234 532574 423854 532658
rect 423234 532338 423266 532574
rect 423502 532338 423586 532574
rect 423822 532338 423854 532574
rect 423234 496894 423854 532338
rect 423234 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 423854 496894
rect 423234 496574 423854 496658
rect 423234 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 423854 496574
rect 423234 460894 423854 496338
rect 423234 460658 423266 460894
rect 423502 460658 423586 460894
rect 423822 460658 423854 460894
rect 423234 460574 423854 460658
rect 423234 460338 423266 460574
rect 423502 460338 423586 460574
rect 423822 460338 423854 460574
rect 423234 442000 423854 460338
rect 426954 680614 427574 711002
rect 444954 710598 445574 711590
rect 444954 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 445574 710598
rect 444954 710278 445574 710362
rect 444954 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 445574 710278
rect 441234 708678 441854 709670
rect 441234 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 441854 708678
rect 441234 708358 441854 708442
rect 441234 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 441854 708358
rect 437514 706758 438134 707750
rect 437514 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 438134 706758
rect 437514 706438 438134 706522
rect 437514 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 438134 706438
rect 426954 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 427574 680614
rect 426954 680294 427574 680378
rect 426954 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 427574 680294
rect 426954 644614 427574 680058
rect 426954 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 427574 644614
rect 426954 644294 427574 644378
rect 426954 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 427574 644294
rect 426954 608614 427574 644058
rect 426954 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 427574 608614
rect 426954 608294 427574 608378
rect 426954 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 427574 608294
rect 426954 572614 427574 608058
rect 426954 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 427574 572614
rect 426954 572294 427574 572378
rect 426954 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 427574 572294
rect 426954 536614 427574 572058
rect 426954 536378 426986 536614
rect 427222 536378 427306 536614
rect 427542 536378 427574 536614
rect 426954 536294 427574 536378
rect 426954 536058 426986 536294
rect 427222 536058 427306 536294
rect 427542 536058 427574 536294
rect 426954 500614 427574 536058
rect 426954 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 427574 500614
rect 426954 500294 427574 500378
rect 426954 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 427574 500294
rect 426954 464614 427574 500058
rect 426954 464378 426986 464614
rect 427222 464378 427306 464614
rect 427542 464378 427574 464614
rect 426954 464294 427574 464378
rect 426954 464058 426986 464294
rect 427222 464058 427306 464294
rect 427542 464058 427574 464294
rect 426954 442000 427574 464058
rect 433794 704838 434414 705830
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 442000 434414 470898
rect 437514 691174 438134 706202
rect 437514 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 438134 691174
rect 437514 690854 438134 690938
rect 437514 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 438134 690854
rect 437514 655174 438134 690618
rect 437514 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 438134 655174
rect 437514 654854 438134 654938
rect 437514 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 438134 654854
rect 437514 619174 438134 654618
rect 437514 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 438134 619174
rect 437514 618854 438134 618938
rect 437514 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 438134 618854
rect 437514 583174 438134 618618
rect 437514 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 438134 583174
rect 437514 582854 438134 582938
rect 437514 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 438134 582854
rect 437514 547174 438134 582618
rect 437514 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 438134 547174
rect 437514 546854 438134 546938
rect 437514 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 438134 546854
rect 437514 511174 438134 546618
rect 437514 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 438134 511174
rect 437514 510854 438134 510938
rect 437514 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 438134 510854
rect 437514 475174 438134 510618
rect 437514 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 438134 475174
rect 437514 474854 438134 474938
rect 437514 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 438134 474854
rect 437514 442000 438134 474618
rect 441234 694894 441854 708122
rect 441234 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 441854 694894
rect 441234 694574 441854 694658
rect 441234 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 441854 694574
rect 441234 658894 441854 694338
rect 441234 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 441854 658894
rect 441234 658574 441854 658658
rect 441234 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 441854 658574
rect 441234 622894 441854 658338
rect 441234 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 441854 622894
rect 441234 622574 441854 622658
rect 441234 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 441854 622574
rect 441234 586894 441854 622338
rect 441234 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 441854 586894
rect 441234 586574 441854 586658
rect 441234 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 441854 586574
rect 441234 550894 441854 586338
rect 441234 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 441854 550894
rect 441234 550574 441854 550658
rect 441234 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 441854 550574
rect 441234 514894 441854 550338
rect 441234 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 441854 514894
rect 441234 514574 441854 514658
rect 441234 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 441854 514574
rect 441234 478894 441854 514338
rect 441234 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 441854 478894
rect 441234 478574 441854 478658
rect 441234 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 441854 478574
rect 441234 442894 441854 478338
rect 441234 442658 441266 442894
rect 441502 442658 441586 442894
rect 441822 442658 441854 442894
rect 441234 442574 441854 442658
rect 441234 442338 441266 442574
rect 441502 442338 441586 442574
rect 441822 442338 441854 442574
rect 441234 442000 441854 442338
rect 444954 698614 445574 710042
rect 462954 711558 463574 711590
rect 462954 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 463574 711558
rect 462954 711238 463574 711322
rect 462954 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 463574 711238
rect 459234 709638 459854 709670
rect 459234 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 459854 709638
rect 459234 709318 459854 709402
rect 459234 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 459854 709318
rect 455514 707718 456134 707750
rect 455514 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 456134 707718
rect 455514 707398 456134 707482
rect 455514 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 456134 707398
rect 444954 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 445574 698614
rect 444954 698294 445574 698378
rect 444954 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 445574 698294
rect 444954 662614 445574 698058
rect 444954 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 445574 662614
rect 444954 662294 445574 662378
rect 444954 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 445574 662294
rect 444954 626614 445574 662058
rect 444954 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 445574 626614
rect 444954 626294 445574 626378
rect 444954 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 445574 626294
rect 444954 590614 445574 626058
rect 444954 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 445574 590614
rect 444954 590294 445574 590378
rect 444954 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 445574 590294
rect 444954 554614 445574 590058
rect 444954 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 445574 554614
rect 444954 554294 445574 554378
rect 444954 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 445574 554294
rect 444954 518614 445574 554058
rect 444954 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 445574 518614
rect 444954 518294 445574 518378
rect 444954 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 445574 518294
rect 444954 482614 445574 518058
rect 444954 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 445574 482614
rect 444954 482294 445574 482378
rect 444954 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 445574 482294
rect 444954 446614 445574 482058
rect 444954 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 445574 446614
rect 444954 446294 445574 446378
rect 444954 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 445574 446294
rect 444954 442000 445574 446058
rect 451794 705798 452414 705830
rect 451794 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 452414 705798
rect 451794 705478 452414 705562
rect 451794 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 452414 705478
rect 451794 669454 452414 705242
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 453454 452414 488898
rect 451794 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 452414 453454
rect 451794 453134 452414 453218
rect 451794 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 452414 453134
rect 451794 442000 452414 452898
rect 455514 673174 456134 707162
rect 455514 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 456134 673174
rect 455514 672854 456134 672938
rect 455514 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 456134 672854
rect 455514 637174 456134 672618
rect 455514 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 456134 637174
rect 455514 636854 456134 636938
rect 455514 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 456134 636854
rect 455514 601174 456134 636618
rect 455514 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 456134 601174
rect 455514 600854 456134 600938
rect 455514 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 456134 600854
rect 455514 565174 456134 600618
rect 455514 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 456134 565174
rect 455514 564854 456134 564938
rect 455514 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 456134 564854
rect 455514 529174 456134 564618
rect 455514 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 456134 529174
rect 455514 528854 456134 528938
rect 455514 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 456134 528854
rect 455514 493174 456134 528618
rect 455514 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 456134 493174
rect 455514 492854 456134 492938
rect 455514 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 456134 492854
rect 455514 457174 456134 492618
rect 455514 456938 455546 457174
rect 455782 456938 455866 457174
rect 456102 456938 456134 457174
rect 455514 456854 456134 456938
rect 455514 456618 455546 456854
rect 455782 456618 455866 456854
rect 456102 456618 456134 456854
rect 455514 442000 456134 456618
rect 459234 676894 459854 709082
rect 459234 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 459854 676894
rect 459234 676574 459854 676658
rect 459234 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 459854 676574
rect 459234 640894 459854 676338
rect 459234 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 459854 640894
rect 459234 640574 459854 640658
rect 459234 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 459854 640574
rect 459234 604894 459854 640338
rect 459234 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 459854 604894
rect 459234 604574 459854 604658
rect 459234 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 459854 604574
rect 459234 568894 459854 604338
rect 459234 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 459854 568894
rect 459234 568574 459854 568658
rect 459234 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 459854 568574
rect 459234 532894 459854 568338
rect 459234 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 459854 532894
rect 459234 532574 459854 532658
rect 459234 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 459854 532574
rect 459234 496894 459854 532338
rect 459234 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 459854 496894
rect 459234 496574 459854 496658
rect 459234 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 459854 496574
rect 459234 460894 459854 496338
rect 459234 460658 459266 460894
rect 459502 460658 459586 460894
rect 459822 460658 459854 460894
rect 459234 460574 459854 460658
rect 459234 460338 459266 460574
rect 459502 460338 459586 460574
rect 459822 460338 459854 460574
rect 459234 442000 459854 460338
rect 462954 680614 463574 711002
rect 480954 710598 481574 711590
rect 480954 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 481574 710598
rect 480954 710278 481574 710362
rect 480954 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 481574 710278
rect 477234 708678 477854 709670
rect 477234 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 477854 708678
rect 477234 708358 477854 708442
rect 477234 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 477854 708358
rect 473514 706758 474134 707750
rect 473514 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 474134 706758
rect 473514 706438 474134 706522
rect 473514 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 474134 706438
rect 462954 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 463574 680614
rect 462954 680294 463574 680378
rect 462954 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 463574 680294
rect 462954 644614 463574 680058
rect 462954 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 463574 644614
rect 462954 644294 463574 644378
rect 462954 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 463574 644294
rect 462954 608614 463574 644058
rect 462954 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 463574 608614
rect 462954 608294 463574 608378
rect 462954 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 463574 608294
rect 462954 572614 463574 608058
rect 462954 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 463574 572614
rect 462954 572294 463574 572378
rect 462954 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 463574 572294
rect 462954 536614 463574 572058
rect 462954 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 463574 536614
rect 462954 536294 463574 536378
rect 462954 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 463574 536294
rect 462954 500614 463574 536058
rect 462954 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 463574 500614
rect 462954 500294 463574 500378
rect 462954 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 463574 500294
rect 462954 464614 463574 500058
rect 462954 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 463574 464614
rect 462954 464294 463574 464378
rect 462954 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 463574 464294
rect 462954 442000 463574 464058
rect 469794 704838 470414 705830
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 442000 470414 470898
rect 473514 691174 474134 706202
rect 473514 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 474134 691174
rect 473514 690854 474134 690938
rect 473514 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 474134 690854
rect 473514 655174 474134 690618
rect 473514 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 474134 655174
rect 473514 654854 474134 654938
rect 473514 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 474134 654854
rect 473514 619174 474134 654618
rect 473514 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 474134 619174
rect 473514 618854 474134 618938
rect 473514 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 474134 618854
rect 473514 583174 474134 618618
rect 473514 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 474134 583174
rect 473514 582854 474134 582938
rect 473514 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 474134 582854
rect 473514 547174 474134 582618
rect 473514 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 474134 547174
rect 473514 546854 474134 546938
rect 473514 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 474134 546854
rect 473514 511174 474134 546618
rect 473514 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 474134 511174
rect 473514 510854 474134 510938
rect 473514 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 474134 510854
rect 473514 475174 474134 510618
rect 473514 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 474134 475174
rect 473514 474854 474134 474938
rect 473514 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 474134 474854
rect 473514 442000 474134 474618
rect 477234 694894 477854 708122
rect 477234 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 477854 694894
rect 477234 694574 477854 694658
rect 477234 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 477854 694574
rect 477234 658894 477854 694338
rect 477234 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 477854 658894
rect 477234 658574 477854 658658
rect 477234 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 477854 658574
rect 477234 622894 477854 658338
rect 477234 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 477854 622894
rect 477234 622574 477854 622658
rect 477234 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 477854 622574
rect 477234 586894 477854 622338
rect 477234 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 477854 586894
rect 477234 586574 477854 586658
rect 477234 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 477854 586574
rect 477234 550894 477854 586338
rect 477234 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 477854 550894
rect 477234 550574 477854 550658
rect 477234 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 477854 550574
rect 477234 514894 477854 550338
rect 477234 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 477854 514894
rect 477234 514574 477854 514658
rect 477234 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 477854 514574
rect 477234 478894 477854 514338
rect 477234 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 477854 478894
rect 477234 478574 477854 478658
rect 477234 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 477854 478574
rect 477234 442894 477854 478338
rect 477234 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 477854 442894
rect 477234 442574 477854 442658
rect 477234 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 477854 442574
rect 477234 442000 477854 442338
rect 480954 698614 481574 710042
rect 498954 711558 499574 711590
rect 498954 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 499574 711558
rect 498954 711238 499574 711322
rect 498954 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 499574 711238
rect 495234 709638 495854 709670
rect 495234 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 495854 709638
rect 495234 709318 495854 709402
rect 495234 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 495854 709318
rect 491514 707718 492134 707750
rect 491514 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 492134 707718
rect 491514 707398 492134 707482
rect 491514 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 492134 707398
rect 480954 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 481574 698614
rect 480954 698294 481574 698378
rect 480954 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 481574 698294
rect 480954 662614 481574 698058
rect 480954 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 481574 662614
rect 480954 662294 481574 662378
rect 480954 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 481574 662294
rect 480954 626614 481574 662058
rect 480954 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 481574 626614
rect 480954 626294 481574 626378
rect 480954 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 481574 626294
rect 480954 590614 481574 626058
rect 480954 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 481574 590614
rect 480954 590294 481574 590378
rect 480954 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 481574 590294
rect 480954 554614 481574 590058
rect 480954 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 481574 554614
rect 480954 554294 481574 554378
rect 480954 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 481574 554294
rect 480954 518614 481574 554058
rect 480954 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 481574 518614
rect 480954 518294 481574 518378
rect 480954 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 481574 518294
rect 480954 482614 481574 518058
rect 480954 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 481574 482614
rect 480954 482294 481574 482378
rect 480954 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 481574 482294
rect 480954 446614 481574 482058
rect 480954 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 481574 446614
rect 480954 446294 481574 446378
rect 480954 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 481574 446294
rect 480954 442000 481574 446058
rect 487794 705798 488414 705830
rect 487794 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 488414 705798
rect 487794 705478 488414 705562
rect 487794 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 488414 705478
rect 487794 669454 488414 705242
rect 491339 700500 491405 700501
rect 491339 700436 491340 700500
rect 491404 700436 491405 700500
rect 491339 700435 491405 700436
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 561454 488414 596898
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 490419 498812 490485 498813
rect 490419 498748 490420 498812
rect 490484 498748 490485 498812
rect 490419 498747 490485 498748
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 453454 488414 488898
rect 487794 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 488414 453454
rect 487794 453134 488414 453218
rect 487794 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 488414 453134
rect 487794 442000 488414 452898
rect 490422 435981 490482 498747
rect 490419 435980 490485 435981
rect 490419 435916 490420 435980
rect 490484 435916 490485 435980
rect 490419 435915 490485 435916
rect 244208 435454 244528 435486
rect 244208 435218 244250 435454
rect 244486 435218 244528 435454
rect 244208 435134 244528 435218
rect 244208 434898 244250 435134
rect 244486 434898 244528 435134
rect 244208 434866 244528 434898
rect 274928 435454 275248 435486
rect 274928 435218 274970 435454
rect 275206 435218 275248 435454
rect 274928 435134 275248 435218
rect 274928 434898 274970 435134
rect 275206 434898 275248 435134
rect 274928 434866 275248 434898
rect 305648 435454 305968 435486
rect 305648 435218 305690 435454
rect 305926 435218 305968 435454
rect 305648 435134 305968 435218
rect 305648 434898 305690 435134
rect 305926 434898 305968 435134
rect 305648 434866 305968 434898
rect 336368 435454 336688 435486
rect 336368 435218 336410 435454
rect 336646 435218 336688 435454
rect 336368 435134 336688 435218
rect 336368 434898 336410 435134
rect 336646 434898 336688 435134
rect 336368 434866 336688 434898
rect 367088 435454 367408 435486
rect 367088 435218 367130 435454
rect 367366 435218 367408 435454
rect 367088 435134 367408 435218
rect 367088 434898 367130 435134
rect 367366 434898 367408 435134
rect 367088 434866 367408 434898
rect 397808 435454 398128 435486
rect 397808 435218 397850 435454
rect 398086 435218 398128 435454
rect 397808 435134 398128 435218
rect 397808 434898 397850 435134
rect 398086 434898 398128 435134
rect 397808 434866 398128 434898
rect 428528 435454 428848 435486
rect 428528 435218 428570 435454
rect 428806 435218 428848 435454
rect 428528 435134 428848 435218
rect 428528 434898 428570 435134
rect 428806 434898 428848 435134
rect 428528 434866 428848 434898
rect 459248 435454 459568 435486
rect 459248 435218 459290 435454
rect 459526 435218 459568 435454
rect 459248 435134 459568 435218
rect 459248 434898 459290 435134
rect 459526 434898 459568 435134
rect 459248 434866 459568 434898
rect 489968 435454 490288 435486
rect 489968 435218 490010 435454
rect 490246 435218 490288 435454
rect 489968 435134 490288 435218
rect 489968 434898 490010 435134
rect 490246 434898 490288 435134
rect 489968 434866 490288 434898
rect 259568 417454 259888 417486
rect 259568 417218 259610 417454
rect 259846 417218 259888 417454
rect 259568 417134 259888 417218
rect 259568 416898 259610 417134
rect 259846 416898 259888 417134
rect 259568 416866 259888 416898
rect 290288 417454 290608 417486
rect 290288 417218 290330 417454
rect 290566 417218 290608 417454
rect 290288 417134 290608 417218
rect 290288 416898 290330 417134
rect 290566 416898 290608 417134
rect 290288 416866 290608 416898
rect 321008 417454 321328 417486
rect 321008 417218 321050 417454
rect 321286 417218 321328 417454
rect 321008 417134 321328 417218
rect 321008 416898 321050 417134
rect 321286 416898 321328 417134
rect 321008 416866 321328 416898
rect 351728 417454 352048 417486
rect 351728 417218 351770 417454
rect 352006 417218 352048 417454
rect 351728 417134 352048 417218
rect 351728 416898 351770 417134
rect 352006 416898 352048 417134
rect 351728 416866 352048 416898
rect 382448 417454 382768 417486
rect 382448 417218 382490 417454
rect 382726 417218 382768 417454
rect 382448 417134 382768 417218
rect 382448 416898 382490 417134
rect 382726 416898 382768 417134
rect 382448 416866 382768 416898
rect 413168 417454 413488 417486
rect 413168 417218 413210 417454
rect 413446 417218 413488 417454
rect 413168 417134 413488 417218
rect 413168 416898 413210 417134
rect 413446 416898 413488 417134
rect 413168 416866 413488 416898
rect 443888 417454 444208 417486
rect 443888 417218 443930 417454
rect 444166 417218 444208 417454
rect 443888 417134 444208 417218
rect 443888 416898 443930 417134
rect 444166 416898 444208 417134
rect 443888 416866 444208 416898
rect 474608 417454 474928 417486
rect 474608 417218 474650 417454
rect 474886 417218 474928 417454
rect 474608 417134 474928 417218
rect 474608 416898 474650 417134
rect 474886 416898 474928 417134
rect 474608 416866 474928 416898
rect 244208 399454 244528 399486
rect 244208 399218 244250 399454
rect 244486 399218 244528 399454
rect 244208 399134 244528 399218
rect 244208 398898 244250 399134
rect 244486 398898 244528 399134
rect 244208 398866 244528 398898
rect 274928 399454 275248 399486
rect 274928 399218 274970 399454
rect 275206 399218 275248 399454
rect 274928 399134 275248 399218
rect 274928 398898 274970 399134
rect 275206 398898 275248 399134
rect 274928 398866 275248 398898
rect 305648 399454 305968 399486
rect 305648 399218 305690 399454
rect 305926 399218 305968 399454
rect 305648 399134 305968 399218
rect 305648 398898 305690 399134
rect 305926 398898 305968 399134
rect 305648 398866 305968 398898
rect 336368 399454 336688 399486
rect 336368 399218 336410 399454
rect 336646 399218 336688 399454
rect 336368 399134 336688 399218
rect 336368 398898 336410 399134
rect 336646 398898 336688 399134
rect 336368 398866 336688 398898
rect 367088 399454 367408 399486
rect 367088 399218 367130 399454
rect 367366 399218 367408 399454
rect 367088 399134 367408 399218
rect 367088 398898 367130 399134
rect 367366 398898 367408 399134
rect 367088 398866 367408 398898
rect 397808 399454 398128 399486
rect 397808 399218 397850 399454
rect 398086 399218 398128 399454
rect 397808 399134 398128 399218
rect 397808 398898 397850 399134
rect 398086 398898 398128 399134
rect 397808 398866 398128 398898
rect 428528 399454 428848 399486
rect 428528 399218 428570 399454
rect 428806 399218 428848 399454
rect 428528 399134 428848 399218
rect 428528 398898 428570 399134
rect 428806 398898 428848 399134
rect 428528 398866 428848 398898
rect 459248 399454 459568 399486
rect 459248 399218 459290 399454
rect 459526 399218 459568 399454
rect 459248 399134 459568 399218
rect 459248 398898 459290 399134
rect 459526 398898 459568 399134
rect 459248 398866 459568 398898
rect 489968 399454 490288 399486
rect 489968 399218 490010 399454
rect 490246 399218 490288 399454
rect 489968 399134 490288 399218
rect 489968 398898 490010 399134
rect 490246 398898 490288 399134
rect 489968 398866 490288 398898
rect 259568 381454 259888 381486
rect 259568 381218 259610 381454
rect 259846 381218 259888 381454
rect 259568 381134 259888 381218
rect 259568 380898 259610 381134
rect 259846 380898 259888 381134
rect 259568 380866 259888 380898
rect 290288 381454 290608 381486
rect 290288 381218 290330 381454
rect 290566 381218 290608 381454
rect 290288 381134 290608 381218
rect 290288 380898 290330 381134
rect 290566 380898 290608 381134
rect 290288 380866 290608 380898
rect 321008 381454 321328 381486
rect 321008 381218 321050 381454
rect 321286 381218 321328 381454
rect 321008 381134 321328 381218
rect 321008 380898 321050 381134
rect 321286 380898 321328 381134
rect 321008 380866 321328 380898
rect 351728 381454 352048 381486
rect 351728 381218 351770 381454
rect 352006 381218 352048 381454
rect 351728 381134 352048 381218
rect 351728 380898 351770 381134
rect 352006 380898 352048 381134
rect 351728 380866 352048 380898
rect 382448 381454 382768 381486
rect 382448 381218 382490 381454
rect 382726 381218 382768 381454
rect 382448 381134 382768 381218
rect 382448 380898 382490 381134
rect 382726 380898 382768 381134
rect 382448 380866 382768 380898
rect 413168 381454 413488 381486
rect 413168 381218 413210 381454
rect 413446 381218 413488 381454
rect 413168 381134 413488 381218
rect 413168 380898 413210 381134
rect 413446 380898 413488 381134
rect 413168 380866 413488 380898
rect 443888 381454 444208 381486
rect 443888 381218 443930 381454
rect 444166 381218 444208 381454
rect 443888 381134 444208 381218
rect 443888 380898 443930 381134
rect 444166 380898 444208 381134
rect 443888 380866 444208 380898
rect 474608 381454 474928 381486
rect 474608 381218 474650 381454
rect 474886 381218 474928 381454
rect 474608 381134 474928 381218
rect 474608 380898 474650 381134
rect 474886 380898 474928 381134
rect 474608 380866 474928 380898
rect 244208 363454 244528 363486
rect 244208 363218 244250 363454
rect 244486 363218 244528 363454
rect 244208 363134 244528 363218
rect 244208 362898 244250 363134
rect 244486 362898 244528 363134
rect 244208 362866 244528 362898
rect 274928 363454 275248 363486
rect 274928 363218 274970 363454
rect 275206 363218 275248 363454
rect 274928 363134 275248 363218
rect 274928 362898 274970 363134
rect 275206 362898 275248 363134
rect 274928 362866 275248 362898
rect 305648 363454 305968 363486
rect 305648 363218 305690 363454
rect 305926 363218 305968 363454
rect 305648 363134 305968 363218
rect 305648 362898 305690 363134
rect 305926 362898 305968 363134
rect 305648 362866 305968 362898
rect 336368 363454 336688 363486
rect 336368 363218 336410 363454
rect 336646 363218 336688 363454
rect 336368 363134 336688 363218
rect 336368 362898 336410 363134
rect 336646 362898 336688 363134
rect 336368 362866 336688 362898
rect 367088 363454 367408 363486
rect 367088 363218 367130 363454
rect 367366 363218 367408 363454
rect 367088 363134 367408 363218
rect 367088 362898 367130 363134
rect 367366 362898 367408 363134
rect 367088 362866 367408 362898
rect 397808 363454 398128 363486
rect 397808 363218 397850 363454
rect 398086 363218 398128 363454
rect 397808 363134 398128 363218
rect 397808 362898 397850 363134
rect 398086 362898 398128 363134
rect 397808 362866 398128 362898
rect 428528 363454 428848 363486
rect 428528 363218 428570 363454
rect 428806 363218 428848 363454
rect 428528 363134 428848 363218
rect 428528 362898 428570 363134
rect 428806 362898 428848 363134
rect 428528 362866 428848 362898
rect 459248 363454 459568 363486
rect 459248 363218 459290 363454
rect 459526 363218 459568 363454
rect 459248 363134 459568 363218
rect 459248 362898 459290 363134
rect 459526 362898 459568 363134
rect 459248 362866 459568 362898
rect 489968 363454 490288 363486
rect 489968 363218 490010 363454
rect 490246 363218 490288 363454
rect 489968 363134 490288 363218
rect 489968 362898 490010 363134
rect 490246 362898 490288 363134
rect 489968 362866 490288 362898
rect 259568 345454 259888 345486
rect 259568 345218 259610 345454
rect 259846 345218 259888 345454
rect 259568 345134 259888 345218
rect 259568 344898 259610 345134
rect 259846 344898 259888 345134
rect 259568 344866 259888 344898
rect 290288 345454 290608 345486
rect 290288 345218 290330 345454
rect 290566 345218 290608 345454
rect 290288 345134 290608 345218
rect 290288 344898 290330 345134
rect 290566 344898 290608 345134
rect 290288 344866 290608 344898
rect 321008 345454 321328 345486
rect 321008 345218 321050 345454
rect 321286 345218 321328 345454
rect 321008 345134 321328 345218
rect 321008 344898 321050 345134
rect 321286 344898 321328 345134
rect 321008 344866 321328 344898
rect 351728 345454 352048 345486
rect 351728 345218 351770 345454
rect 352006 345218 352048 345454
rect 351728 345134 352048 345218
rect 351728 344898 351770 345134
rect 352006 344898 352048 345134
rect 351728 344866 352048 344898
rect 382448 345454 382768 345486
rect 382448 345218 382490 345454
rect 382726 345218 382768 345454
rect 382448 345134 382768 345218
rect 382448 344898 382490 345134
rect 382726 344898 382768 345134
rect 382448 344866 382768 344898
rect 413168 345454 413488 345486
rect 413168 345218 413210 345454
rect 413446 345218 413488 345454
rect 413168 345134 413488 345218
rect 413168 344898 413210 345134
rect 413446 344898 413488 345134
rect 413168 344866 413488 344898
rect 443888 345454 444208 345486
rect 443888 345218 443930 345454
rect 444166 345218 444208 345454
rect 443888 345134 444208 345218
rect 443888 344898 443930 345134
rect 444166 344898 444208 345134
rect 443888 344866 444208 344898
rect 474608 345454 474928 345486
rect 474608 345218 474650 345454
rect 474886 345218 474928 345454
rect 474608 345134 474928 345218
rect 474608 344898 474650 345134
rect 474886 344898 474928 345134
rect 474608 344866 474928 344898
rect 244208 327454 244528 327486
rect 244208 327218 244250 327454
rect 244486 327218 244528 327454
rect 244208 327134 244528 327218
rect 244208 326898 244250 327134
rect 244486 326898 244528 327134
rect 244208 326866 244528 326898
rect 274928 327454 275248 327486
rect 274928 327218 274970 327454
rect 275206 327218 275248 327454
rect 274928 327134 275248 327218
rect 274928 326898 274970 327134
rect 275206 326898 275248 327134
rect 274928 326866 275248 326898
rect 305648 327454 305968 327486
rect 305648 327218 305690 327454
rect 305926 327218 305968 327454
rect 305648 327134 305968 327218
rect 305648 326898 305690 327134
rect 305926 326898 305968 327134
rect 305648 326866 305968 326898
rect 336368 327454 336688 327486
rect 336368 327218 336410 327454
rect 336646 327218 336688 327454
rect 336368 327134 336688 327218
rect 336368 326898 336410 327134
rect 336646 326898 336688 327134
rect 336368 326866 336688 326898
rect 367088 327454 367408 327486
rect 367088 327218 367130 327454
rect 367366 327218 367408 327454
rect 367088 327134 367408 327218
rect 367088 326898 367130 327134
rect 367366 326898 367408 327134
rect 367088 326866 367408 326898
rect 397808 327454 398128 327486
rect 397808 327218 397850 327454
rect 398086 327218 398128 327454
rect 397808 327134 398128 327218
rect 397808 326898 397850 327134
rect 398086 326898 398128 327134
rect 397808 326866 398128 326898
rect 428528 327454 428848 327486
rect 428528 327218 428570 327454
rect 428806 327218 428848 327454
rect 428528 327134 428848 327218
rect 428528 326898 428570 327134
rect 428806 326898 428848 327134
rect 428528 326866 428848 326898
rect 459248 327454 459568 327486
rect 459248 327218 459290 327454
rect 459526 327218 459568 327454
rect 459248 327134 459568 327218
rect 459248 326898 459290 327134
rect 459526 326898 459568 327134
rect 459248 326866 459568 326898
rect 489968 327454 490288 327486
rect 489968 327218 490010 327454
rect 490246 327218 490288 327454
rect 489968 327134 490288 327218
rect 489968 326898 490010 327134
rect 490246 326898 490288 327134
rect 489968 326866 490288 326898
rect 259568 309454 259888 309486
rect 259568 309218 259610 309454
rect 259846 309218 259888 309454
rect 259568 309134 259888 309218
rect 259568 308898 259610 309134
rect 259846 308898 259888 309134
rect 259568 308866 259888 308898
rect 290288 309454 290608 309486
rect 290288 309218 290330 309454
rect 290566 309218 290608 309454
rect 290288 309134 290608 309218
rect 290288 308898 290330 309134
rect 290566 308898 290608 309134
rect 290288 308866 290608 308898
rect 321008 309454 321328 309486
rect 321008 309218 321050 309454
rect 321286 309218 321328 309454
rect 321008 309134 321328 309218
rect 321008 308898 321050 309134
rect 321286 308898 321328 309134
rect 321008 308866 321328 308898
rect 351728 309454 352048 309486
rect 351728 309218 351770 309454
rect 352006 309218 352048 309454
rect 351728 309134 352048 309218
rect 351728 308898 351770 309134
rect 352006 308898 352048 309134
rect 351728 308866 352048 308898
rect 382448 309454 382768 309486
rect 382448 309218 382490 309454
rect 382726 309218 382768 309454
rect 382448 309134 382768 309218
rect 382448 308898 382490 309134
rect 382726 308898 382768 309134
rect 382448 308866 382768 308898
rect 413168 309454 413488 309486
rect 413168 309218 413210 309454
rect 413446 309218 413488 309454
rect 413168 309134 413488 309218
rect 413168 308898 413210 309134
rect 413446 308898 413488 309134
rect 413168 308866 413488 308898
rect 443888 309454 444208 309486
rect 443888 309218 443930 309454
rect 444166 309218 444208 309454
rect 443888 309134 444208 309218
rect 443888 308898 443930 309134
rect 444166 308898 444208 309134
rect 443888 308866 444208 308898
rect 474608 309454 474928 309486
rect 474608 309218 474650 309454
rect 474886 309218 474928 309454
rect 474608 309134 474928 309218
rect 474608 308898 474650 309134
rect 474886 308898 474928 309134
rect 474608 308866 474928 308898
rect 244208 291454 244528 291486
rect 244208 291218 244250 291454
rect 244486 291218 244528 291454
rect 244208 291134 244528 291218
rect 244208 290898 244250 291134
rect 244486 290898 244528 291134
rect 244208 290866 244528 290898
rect 274928 291454 275248 291486
rect 274928 291218 274970 291454
rect 275206 291218 275248 291454
rect 274928 291134 275248 291218
rect 274928 290898 274970 291134
rect 275206 290898 275248 291134
rect 274928 290866 275248 290898
rect 305648 291454 305968 291486
rect 305648 291218 305690 291454
rect 305926 291218 305968 291454
rect 305648 291134 305968 291218
rect 305648 290898 305690 291134
rect 305926 290898 305968 291134
rect 305648 290866 305968 290898
rect 336368 291454 336688 291486
rect 336368 291218 336410 291454
rect 336646 291218 336688 291454
rect 336368 291134 336688 291218
rect 336368 290898 336410 291134
rect 336646 290898 336688 291134
rect 336368 290866 336688 290898
rect 367088 291454 367408 291486
rect 367088 291218 367130 291454
rect 367366 291218 367408 291454
rect 367088 291134 367408 291218
rect 367088 290898 367130 291134
rect 367366 290898 367408 291134
rect 367088 290866 367408 290898
rect 397808 291454 398128 291486
rect 397808 291218 397850 291454
rect 398086 291218 398128 291454
rect 397808 291134 398128 291218
rect 397808 290898 397850 291134
rect 398086 290898 398128 291134
rect 397808 290866 398128 290898
rect 428528 291454 428848 291486
rect 428528 291218 428570 291454
rect 428806 291218 428848 291454
rect 428528 291134 428848 291218
rect 428528 290898 428570 291134
rect 428806 290898 428848 291134
rect 428528 290866 428848 290898
rect 459248 291454 459568 291486
rect 459248 291218 459290 291454
rect 459526 291218 459568 291454
rect 459248 291134 459568 291218
rect 459248 290898 459290 291134
rect 459526 290898 459568 291134
rect 459248 290866 459568 290898
rect 489968 291454 490288 291486
rect 489968 291218 490010 291454
rect 490246 291218 490288 291454
rect 489968 291134 490288 291218
rect 489968 290898 490010 291134
rect 490246 290898 490288 291134
rect 489968 290866 490288 290898
rect 259568 273454 259888 273486
rect 259568 273218 259610 273454
rect 259846 273218 259888 273454
rect 259568 273134 259888 273218
rect 259568 272898 259610 273134
rect 259846 272898 259888 273134
rect 259568 272866 259888 272898
rect 290288 273454 290608 273486
rect 290288 273218 290330 273454
rect 290566 273218 290608 273454
rect 290288 273134 290608 273218
rect 290288 272898 290330 273134
rect 290566 272898 290608 273134
rect 290288 272866 290608 272898
rect 321008 273454 321328 273486
rect 321008 273218 321050 273454
rect 321286 273218 321328 273454
rect 321008 273134 321328 273218
rect 321008 272898 321050 273134
rect 321286 272898 321328 273134
rect 321008 272866 321328 272898
rect 351728 273454 352048 273486
rect 351728 273218 351770 273454
rect 352006 273218 352048 273454
rect 351728 273134 352048 273218
rect 351728 272898 351770 273134
rect 352006 272898 352048 273134
rect 351728 272866 352048 272898
rect 382448 273454 382768 273486
rect 382448 273218 382490 273454
rect 382726 273218 382768 273454
rect 382448 273134 382768 273218
rect 382448 272898 382490 273134
rect 382726 272898 382768 273134
rect 382448 272866 382768 272898
rect 413168 273454 413488 273486
rect 413168 273218 413210 273454
rect 413446 273218 413488 273454
rect 413168 273134 413488 273218
rect 413168 272898 413210 273134
rect 413446 272898 413488 273134
rect 413168 272866 413488 272898
rect 443888 273454 444208 273486
rect 443888 273218 443930 273454
rect 444166 273218 444208 273454
rect 443888 273134 444208 273218
rect 443888 272898 443930 273134
rect 444166 272898 444208 273134
rect 443888 272866 444208 272898
rect 474608 273454 474928 273486
rect 474608 273218 474650 273454
rect 474886 273218 474928 273454
rect 474608 273134 474928 273218
rect 474608 272898 474650 273134
rect 474886 272898 474928 273134
rect 474608 272866 474928 272898
rect 244208 255454 244528 255486
rect 244208 255218 244250 255454
rect 244486 255218 244528 255454
rect 244208 255134 244528 255218
rect 244208 254898 244250 255134
rect 244486 254898 244528 255134
rect 244208 254866 244528 254898
rect 274928 255454 275248 255486
rect 274928 255218 274970 255454
rect 275206 255218 275248 255454
rect 274928 255134 275248 255218
rect 274928 254898 274970 255134
rect 275206 254898 275248 255134
rect 274928 254866 275248 254898
rect 305648 255454 305968 255486
rect 305648 255218 305690 255454
rect 305926 255218 305968 255454
rect 305648 255134 305968 255218
rect 305648 254898 305690 255134
rect 305926 254898 305968 255134
rect 305648 254866 305968 254898
rect 336368 255454 336688 255486
rect 336368 255218 336410 255454
rect 336646 255218 336688 255454
rect 336368 255134 336688 255218
rect 336368 254898 336410 255134
rect 336646 254898 336688 255134
rect 336368 254866 336688 254898
rect 367088 255454 367408 255486
rect 367088 255218 367130 255454
rect 367366 255218 367408 255454
rect 367088 255134 367408 255218
rect 367088 254898 367130 255134
rect 367366 254898 367408 255134
rect 367088 254866 367408 254898
rect 397808 255454 398128 255486
rect 397808 255218 397850 255454
rect 398086 255218 398128 255454
rect 397808 255134 398128 255218
rect 397808 254898 397850 255134
rect 398086 254898 398128 255134
rect 397808 254866 398128 254898
rect 428528 255454 428848 255486
rect 428528 255218 428570 255454
rect 428806 255218 428848 255454
rect 428528 255134 428848 255218
rect 428528 254898 428570 255134
rect 428806 254898 428848 255134
rect 428528 254866 428848 254898
rect 459248 255454 459568 255486
rect 459248 255218 459290 255454
rect 459526 255218 459568 255454
rect 459248 255134 459568 255218
rect 459248 254898 459290 255134
rect 459526 254898 459568 255134
rect 459248 254866 459568 254898
rect 489968 255454 490288 255486
rect 489968 255218 490010 255454
rect 490246 255218 490288 255454
rect 489968 255134 490288 255218
rect 489968 254898 490010 255134
rect 490246 254898 490288 255134
rect 489968 254866 490288 254898
rect 259568 237454 259888 237486
rect 259568 237218 259610 237454
rect 259846 237218 259888 237454
rect 259568 237134 259888 237218
rect 259568 236898 259610 237134
rect 259846 236898 259888 237134
rect 259568 236866 259888 236898
rect 290288 237454 290608 237486
rect 290288 237218 290330 237454
rect 290566 237218 290608 237454
rect 290288 237134 290608 237218
rect 290288 236898 290330 237134
rect 290566 236898 290608 237134
rect 290288 236866 290608 236898
rect 321008 237454 321328 237486
rect 321008 237218 321050 237454
rect 321286 237218 321328 237454
rect 321008 237134 321328 237218
rect 321008 236898 321050 237134
rect 321286 236898 321328 237134
rect 321008 236866 321328 236898
rect 351728 237454 352048 237486
rect 351728 237218 351770 237454
rect 352006 237218 352048 237454
rect 351728 237134 352048 237218
rect 351728 236898 351770 237134
rect 352006 236898 352048 237134
rect 351728 236866 352048 236898
rect 382448 237454 382768 237486
rect 382448 237218 382490 237454
rect 382726 237218 382768 237454
rect 382448 237134 382768 237218
rect 382448 236898 382490 237134
rect 382726 236898 382768 237134
rect 382448 236866 382768 236898
rect 413168 237454 413488 237486
rect 413168 237218 413210 237454
rect 413446 237218 413488 237454
rect 413168 237134 413488 237218
rect 413168 236898 413210 237134
rect 413446 236898 413488 237134
rect 413168 236866 413488 236898
rect 443888 237454 444208 237486
rect 443888 237218 443930 237454
rect 444166 237218 444208 237454
rect 443888 237134 444208 237218
rect 443888 236898 443930 237134
rect 444166 236898 444208 237134
rect 443888 236866 444208 236898
rect 474608 237454 474928 237486
rect 474608 237218 474650 237454
rect 474886 237218 474928 237454
rect 474608 237134 474928 237218
rect 474608 236898 474650 237134
rect 474886 236898 474928 237134
rect 474608 236866 474928 236898
rect 244208 219454 244528 219486
rect 244208 219218 244250 219454
rect 244486 219218 244528 219454
rect 244208 219134 244528 219218
rect 244208 218898 244250 219134
rect 244486 218898 244528 219134
rect 244208 218866 244528 218898
rect 274928 219454 275248 219486
rect 274928 219218 274970 219454
rect 275206 219218 275248 219454
rect 274928 219134 275248 219218
rect 274928 218898 274970 219134
rect 275206 218898 275248 219134
rect 274928 218866 275248 218898
rect 305648 219454 305968 219486
rect 305648 219218 305690 219454
rect 305926 219218 305968 219454
rect 305648 219134 305968 219218
rect 305648 218898 305690 219134
rect 305926 218898 305968 219134
rect 305648 218866 305968 218898
rect 336368 219454 336688 219486
rect 336368 219218 336410 219454
rect 336646 219218 336688 219454
rect 336368 219134 336688 219218
rect 336368 218898 336410 219134
rect 336646 218898 336688 219134
rect 336368 218866 336688 218898
rect 367088 219454 367408 219486
rect 367088 219218 367130 219454
rect 367366 219218 367408 219454
rect 367088 219134 367408 219218
rect 367088 218898 367130 219134
rect 367366 218898 367408 219134
rect 367088 218866 367408 218898
rect 397808 219454 398128 219486
rect 397808 219218 397850 219454
rect 398086 219218 398128 219454
rect 397808 219134 398128 219218
rect 397808 218898 397850 219134
rect 398086 218898 398128 219134
rect 397808 218866 398128 218898
rect 428528 219454 428848 219486
rect 428528 219218 428570 219454
rect 428806 219218 428848 219454
rect 428528 219134 428848 219218
rect 428528 218898 428570 219134
rect 428806 218898 428848 219134
rect 428528 218866 428848 218898
rect 459248 219454 459568 219486
rect 459248 219218 459290 219454
rect 459526 219218 459568 219454
rect 459248 219134 459568 219218
rect 459248 218898 459290 219134
rect 459526 218898 459568 219134
rect 459248 218866 459568 218898
rect 489968 219454 490288 219486
rect 489968 219218 490010 219454
rect 490246 219218 490288 219454
rect 489968 219134 490288 219218
rect 489968 218898 490010 219134
rect 490246 218898 490288 219134
rect 489968 218866 490288 218898
rect 259568 201454 259888 201486
rect 259568 201218 259610 201454
rect 259846 201218 259888 201454
rect 259568 201134 259888 201218
rect 259568 200898 259610 201134
rect 259846 200898 259888 201134
rect 259568 200866 259888 200898
rect 290288 201454 290608 201486
rect 290288 201218 290330 201454
rect 290566 201218 290608 201454
rect 290288 201134 290608 201218
rect 290288 200898 290330 201134
rect 290566 200898 290608 201134
rect 290288 200866 290608 200898
rect 321008 201454 321328 201486
rect 321008 201218 321050 201454
rect 321286 201218 321328 201454
rect 321008 201134 321328 201218
rect 321008 200898 321050 201134
rect 321286 200898 321328 201134
rect 321008 200866 321328 200898
rect 351728 201454 352048 201486
rect 351728 201218 351770 201454
rect 352006 201218 352048 201454
rect 351728 201134 352048 201218
rect 351728 200898 351770 201134
rect 352006 200898 352048 201134
rect 351728 200866 352048 200898
rect 382448 201454 382768 201486
rect 382448 201218 382490 201454
rect 382726 201218 382768 201454
rect 382448 201134 382768 201218
rect 382448 200898 382490 201134
rect 382726 200898 382768 201134
rect 382448 200866 382768 200898
rect 413168 201454 413488 201486
rect 413168 201218 413210 201454
rect 413446 201218 413488 201454
rect 413168 201134 413488 201218
rect 413168 200898 413210 201134
rect 413446 200898 413488 201134
rect 413168 200866 413488 200898
rect 443888 201454 444208 201486
rect 443888 201218 443930 201454
rect 444166 201218 444208 201454
rect 443888 201134 444208 201218
rect 443888 200898 443930 201134
rect 444166 200898 444208 201134
rect 443888 200866 444208 200898
rect 474608 201454 474928 201486
rect 474608 201218 474650 201454
rect 474886 201218 474928 201454
rect 474608 201134 474928 201218
rect 474608 200898 474650 201134
rect 474886 200898 474928 201134
rect 474608 200866 474928 200898
rect 244208 183454 244528 183486
rect 244208 183218 244250 183454
rect 244486 183218 244528 183454
rect 244208 183134 244528 183218
rect 244208 182898 244250 183134
rect 244486 182898 244528 183134
rect 244208 182866 244528 182898
rect 274928 183454 275248 183486
rect 274928 183218 274970 183454
rect 275206 183218 275248 183454
rect 274928 183134 275248 183218
rect 274928 182898 274970 183134
rect 275206 182898 275248 183134
rect 274928 182866 275248 182898
rect 305648 183454 305968 183486
rect 305648 183218 305690 183454
rect 305926 183218 305968 183454
rect 305648 183134 305968 183218
rect 305648 182898 305690 183134
rect 305926 182898 305968 183134
rect 305648 182866 305968 182898
rect 336368 183454 336688 183486
rect 336368 183218 336410 183454
rect 336646 183218 336688 183454
rect 336368 183134 336688 183218
rect 336368 182898 336410 183134
rect 336646 182898 336688 183134
rect 336368 182866 336688 182898
rect 367088 183454 367408 183486
rect 367088 183218 367130 183454
rect 367366 183218 367408 183454
rect 367088 183134 367408 183218
rect 367088 182898 367130 183134
rect 367366 182898 367408 183134
rect 367088 182866 367408 182898
rect 397808 183454 398128 183486
rect 397808 183218 397850 183454
rect 398086 183218 398128 183454
rect 397808 183134 398128 183218
rect 397808 182898 397850 183134
rect 398086 182898 398128 183134
rect 397808 182866 398128 182898
rect 428528 183454 428848 183486
rect 428528 183218 428570 183454
rect 428806 183218 428848 183454
rect 428528 183134 428848 183218
rect 428528 182898 428570 183134
rect 428806 182898 428848 183134
rect 428528 182866 428848 182898
rect 459248 183454 459568 183486
rect 459248 183218 459290 183454
rect 459526 183218 459568 183454
rect 459248 183134 459568 183218
rect 459248 182898 459290 183134
rect 459526 182898 459568 183134
rect 459248 182866 459568 182898
rect 489968 183454 490288 183486
rect 489968 183218 490010 183454
rect 490246 183218 490288 183454
rect 489968 183134 490288 183218
rect 489968 182898 490010 183134
rect 490246 182898 490288 183134
rect 489968 182866 490288 182898
rect 490419 182068 490485 182069
rect 490419 182004 490420 182068
rect 490484 182004 490485 182068
rect 490419 182003 490485 182004
rect 239259 179076 239325 179077
rect 239259 179012 239260 179076
rect 239324 179012 239325 179076
rect 239259 179011 239325 179012
rect 490422 178941 490482 182003
rect 490419 178940 490485 178941
rect 490419 178876 490420 178940
rect 490484 178876 490485 178940
rect 490419 178875 490485 178876
rect 491342 178805 491402 700435
rect 491514 673174 492134 707162
rect 492811 700364 492877 700365
rect 492811 700300 492812 700364
rect 492876 700300 492877 700364
rect 492811 700299 492877 700300
rect 491514 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 492134 673174
rect 491514 672854 492134 672938
rect 491514 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 492134 672854
rect 491514 637174 492134 672618
rect 491514 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 492134 637174
rect 491514 636854 492134 636938
rect 491514 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 492134 636854
rect 491514 601174 492134 636618
rect 491514 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 492134 601174
rect 491514 600854 492134 600938
rect 491514 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 492134 600854
rect 491514 565174 492134 600618
rect 491514 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 492134 565174
rect 491514 564854 492134 564938
rect 491514 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 492134 564854
rect 491514 529174 492134 564618
rect 491514 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 492134 529174
rect 491514 528854 492134 528938
rect 491514 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 492134 528854
rect 491514 493174 492134 528618
rect 491514 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 492134 493174
rect 491514 492854 492134 492938
rect 491514 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 492134 492854
rect 491514 457174 492134 492618
rect 491514 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 492134 457174
rect 491514 456854 492134 456938
rect 491514 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 492134 456854
rect 491514 442000 492134 456618
rect 491523 435980 491589 435981
rect 491523 435916 491524 435980
rect 491588 435916 491589 435980
rect 491523 435915 491589 435916
rect 491526 182069 491586 435915
rect 491523 182068 491589 182069
rect 491523 182004 491524 182068
rect 491588 182004 491589 182068
rect 491523 182003 491589 182004
rect 491339 178804 491405 178805
rect 491339 178740 491340 178804
rect 491404 178740 491405 178804
rect 491339 178739 491405 178740
rect 492814 178669 492874 700299
rect 495234 676894 495854 709082
rect 495234 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 495854 676894
rect 495234 676574 495854 676658
rect 495234 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 495854 676574
rect 495234 640894 495854 676338
rect 495234 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 495854 640894
rect 495234 640574 495854 640658
rect 495234 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 495854 640574
rect 495234 604894 495854 640338
rect 495234 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 495854 604894
rect 495234 604574 495854 604658
rect 495234 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 495854 604574
rect 495234 568894 495854 604338
rect 495234 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 495854 568894
rect 495234 568574 495854 568658
rect 495234 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 495854 568574
rect 495234 532894 495854 568338
rect 495234 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 495854 532894
rect 495234 532574 495854 532658
rect 495234 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 495854 532574
rect 495234 496894 495854 532338
rect 495234 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 495854 496894
rect 495234 496574 495854 496658
rect 495234 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 495854 496574
rect 494099 488612 494165 488613
rect 494099 488548 494100 488612
rect 494164 488548 494165 488612
rect 494099 488547 494165 488548
rect 494102 179485 494162 488547
rect 495234 460894 495854 496338
rect 495234 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 495854 460894
rect 495234 460574 495854 460658
rect 495234 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 495854 460574
rect 495234 442000 495854 460338
rect 498954 680614 499574 711002
rect 516954 710598 517574 711590
rect 516954 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 517574 710598
rect 516954 710278 517574 710362
rect 516954 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 517574 710278
rect 513234 708678 513854 709670
rect 513234 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 513854 708678
rect 513234 708358 513854 708442
rect 513234 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 513854 708358
rect 509514 706758 510134 707750
rect 509514 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 510134 706758
rect 509514 706438 510134 706522
rect 509514 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 510134 706438
rect 498954 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 499574 680614
rect 498954 680294 499574 680378
rect 498954 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 499574 680294
rect 498954 644614 499574 680058
rect 498954 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 499574 644614
rect 498954 644294 499574 644378
rect 498954 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 499574 644294
rect 498954 608614 499574 644058
rect 498954 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 499574 608614
rect 498954 608294 499574 608378
rect 498954 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 499574 608294
rect 498954 572614 499574 608058
rect 498954 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 499574 572614
rect 498954 572294 499574 572378
rect 498954 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 499574 572294
rect 498954 536614 499574 572058
rect 498954 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 499574 536614
rect 498954 536294 499574 536378
rect 498954 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 499574 536294
rect 498954 500614 499574 536058
rect 498954 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 499574 500614
rect 498954 500294 499574 500378
rect 498954 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 499574 500294
rect 498954 464614 499574 500058
rect 498954 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 499574 464614
rect 498954 464294 499574 464378
rect 498954 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 499574 464294
rect 498954 442000 499574 464058
rect 505794 704838 506414 705830
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 494099 179484 494165 179485
rect 494099 179420 494100 179484
rect 494164 179420 494165 179484
rect 494099 179419 494165 179420
rect 492811 178668 492877 178669
rect 492811 178604 492812 178668
rect 492876 178604 492877 178668
rect 492811 178603 492877 178604
rect 235794 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 236414 165454
rect 235794 165134 236414 165218
rect 235794 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 236414 165134
rect 235794 129454 236414 164898
rect 235794 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 236414 129454
rect 235794 129134 236414 129218
rect 235794 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 236414 129134
rect 235794 93454 236414 128898
rect 235794 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 236414 93454
rect 235794 93134 236414 93218
rect 235794 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 236414 93134
rect 235794 57454 236414 92898
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -1306 236414 20898
rect 235794 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 236414 -1306
rect 235794 -1626 236414 -1542
rect 235794 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 236414 -1626
rect 235794 -1894 236414 -1862
rect 239514 169174 240134 178000
rect 239514 168938 239546 169174
rect 239782 168938 239866 169174
rect 240102 168938 240134 169174
rect 239514 168854 240134 168938
rect 239514 168618 239546 168854
rect 239782 168618 239866 168854
rect 240102 168618 240134 168854
rect 239514 133174 240134 168618
rect 239514 132938 239546 133174
rect 239782 132938 239866 133174
rect 240102 132938 240134 133174
rect 239514 132854 240134 132938
rect 239514 132618 239546 132854
rect 239782 132618 239866 132854
rect 240102 132618 240134 132854
rect 239514 97174 240134 132618
rect 239514 96938 239546 97174
rect 239782 96938 239866 97174
rect 240102 96938 240134 97174
rect 239514 96854 240134 96938
rect 239514 96618 239546 96854
rect 239782 96618 239866 96854
rect 240102 96618 240134 96854
rect 239514 61174 240134 96618
rect 239514 60938 239546 61174
rect 239782 60938 239866 61174
rect 240102 60938 240134 61174
rect 239514 60854 240134 60938
rect 239514 60618 239546 60854
rect 239782 60618 239866 60854
rect 240102 60618 240134 60854
rect 239514 25174 240134 60618
rect 239514 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 240134 25174
rect 239514 24854 240134 24938
rect 239514 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 240134 24854
rect 239514 -3226 240134 24618
rect 239514 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 240134 -3226
rect 239514 -3546 240134 -3462
rect 239514 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 240134 -3546
rect 239514 -3814 240134 -3782
rect 243234 172894 243854 178000
rect 243234 172658 243266 172894
rect 243502 172658 243586 172894
rect 243822 172658 243854 172894
rect 243234 172574 243854 172658
rect 243234 172338 243266 172574
rect 243502 172338 243586 172574
rect 243822 172338 243854 172574
rect 243234 136894 243854 172338
rect 243234 136658 243266 136894
rect 243502 136658 243586 136894
rect 243822 136658 243854 136894
rect 243234 136574 243854 136658
rect 243234 136338 243266 136574
rect 243502 136338 243586 136574
rect 243822 136338 243854 136574
rect 243234 100894 243854 136338
rect 243234 100658 243266 100894
rect 243502 100658 243586 100894
rect 243822 100658 243854 100894
rect 243234 100574 243854 100658
rect 243234 100338 243266 100574
rect 243502 100338 243586 100574
rect 243822 100338 243854 100574
rect 243234 64894 243854 100338
rect 243234 64658 243266 64894
rect 243502 64658 243586 64894
rect 243822 64658 243854 64894
rect 243234 64574 243854 64658
rect 243234 64338 243266 64574
rect 243502 64338 243586 64574
rect 243822 64338 243854 64574
rect 243234 28894 243854 64338
rect 243234 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 243854 28894
rect 243234 28574 243854 28658
rect 243234 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 243854 28574
rect 243234 -5146 243854 28338
rect 243234 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 243854 -5146
rect 243234 -5466 243854 -5382
rect 243234 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 243854 -5466
rect 243234 -5734 243854 -5702
rect 246954 176614 247574 178000
rect 246954 176378 246986 176614
rect 247222 176378 247306 176614
rect 247542 176378 247574 176614
rect 246954 176294 247574 176378
rect 246954 176058 246986 176294
rect 247222 176058 247306 176294
rect 247542 176058 247574 176294
rect 246954 140614 247574 176058
rect 246954 140378 246986 140614
rect 247222 140378 247306 140614
rect 247542 140378 247574 140614
rect 246954 140294 247574 140378
rect 246954 140058 246986 140294
rect 247222 140058 247306 140294
rect 247542 140058 247574 140294
rect 246954 104614 247574 140058
rect 246954 104378 246986 104614
rect 247222 104378 247306 104614
rect 247542 104378 247574 104614
rect 246954 104294 247574 104378
rect 246954 104058 246986 104294
rect 247222 104058 247306 104294
rect 247542 104058 247574 104294
rect 246954 68614 247574 104058
rect 246954 68378 246986 68614
rect 247222 68378 247306 68614
rect 247542 68378 247574 68614
rect 246954 68294 247574 68378
rect 246954 68058 246986 68294
rect 247222 68058 247306 68294
rect 247542 68058 247574 68294
rect 246954 32614 247574 68058
rect 246954 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 247574 32614
rect 246954 32294 247574 32378
rect 246954 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 247574 32294
rect 228954 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 229574 -6106
rect 228954 -6426 229574 -6342
rect 228954 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 229574 -6426
rect 228954 -7654 229574 -6662
rect 246954 -7066 247574 32058
rect 253794 147454 254414 178000
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 253794 111454 254414 146898
rect 253794 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 254414 111454
rect 253794 111134 254414 111218
rect 253794 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 254414 111134
rect 253794 75454 254414 110898
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -1894 254414 -902
rect 257514 151174 258134 178000
rect 257514 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 258134 151174
rect 257514 150854 258134 150938
rect 257514 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 258134 150854
rect 257514 115174 258134 150618
rect 257514 114938 257546 115174
rect 257782 114938 257866 115174
rect 258102 114938 258134 115174
rect 257514 114854 258134 114938
rect 257514 114618 257546 114854
rect 257782 114618 257866 114854
rect 258102 114618 258134 114854
rect 257514 79174 258134 114618
rect 257514 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 258134 79174
rect 257514 78854 258134 78938
rect 257514 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 258134 78854
rect 257514 43174 258134 78618
rect 257514 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 258134 43174
rect 257514 42854 258134 42938
rect 257514 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 258134 42854
rect 257514 7174 258134 42618
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 257514 -2266 258134 6618
rect 257514 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 258134 -2266
rect 257514 -2586 258134 -2502
rect 257514 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 258134 -2586
rect 257514 -3814 258134 -2822
rect 261234 154894 261854 178000
rect 261234 154658 261266 154894
rect 261502 154658 261586 154894
rect 261822 154658 261854 154894
rect 261234 154574 261854 154658
rect 261234 154338 261266 154574
rect 261502 154338 261586 154574
rect 261822 154338 261854 154574
rect 261234 118894 261854 154338
rect 261234 118658 261266 118894
rect 261502 118658 261586 118894
rect 261822 118658 261854 118894
rect 261234 118574 261854 118658
rect 261234 118338 261266 118574
rect 261502 118338 261586 118574
rect 261822 118338 261854 118574
rect 261234 82894 261854 118338
rect 261234 82658 261266 82894
rect 261502 82658 261586 82894
rect 261822 82658 261854 82894
rect 261234 82574 261854 82658
rect 261234 82338 261266 82574
rect 261502 82338 261586 82574
rect 261822 82338 261854 82574
rect 261234 46894 261854 82338
rect 261234 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 261854 46894
rect 261234 46574 261854 46658
rect 261234 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 261854 46574
rect 261234 10894 261854 46338
rect 261234 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 261854 10894
rect 261234 10574 261854 10658
rect 261234 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 261854 10574
rect 261234 -4186 261854 10338
rect 261234 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 261854 -4186
rect 261234 -4506 261854 -4422
rect 261234 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 261854 -4506
rect 261234 -5734 261854 -4742
rect 264954 158614 265574 178000
rect 264954 158378 264986 158614
rect 265222 158378 265306 158614
rect 265542 158378 265574 158614
rect 264954 158294 265574 158378
rect 264954 158058 264986 158294
rect 265222 158058 265306 158294
rect 265542 158058 265574 158294
rect 264954 122614 265574 158058
rect 264954 122378 264986 122614
rect 265222 122378 265306 122614
rect 265542 122378 265574 122614
rect 264954 122294 265574 122378
rect 264954 122058 264986 122294
rect 265222 122058 265306 122294
rect 265542 122058 265574 122294
rect 264954 86614 265574 122058
rect 264954 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 265574 86614
rect 264954 86294 265574 86378
rect 264954 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 265574 86294
rect 264954 50614 265574 86058
rect 264954 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 265574 50614
rect 264954 50294 265574 50378
rect 264954 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 265574 50294
rect 264954 14614 265574 50058
rect 264954 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 265574 14614
rect 264954 14294 265574 14378
rect 264954 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 265574 14294
rect 246954 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 247574 -7066
rect 246954 -7386 247574 -7302
rect 246954 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 247574 -7386
rect 246954 -7654 247574 -7622
rect 264954 -6106 265574 14058
rect 271794 165454 272414 178000
rect 271794 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 272414 165454
rect 271794 165134 272414 165218
rect 271794 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 272414 165134
rect 271794 129454 272414 164898
rect 271794 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 272414 129454
rect 271794 129134 272414 129218
rect 271794 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 272414 129134
rect 271794 93454 272414 128898
rect 271794 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 272414 93454
rect 271794 93134 272414 93218
rect 271794 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 272414 93134
rect 271794 57454 272414 92898
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -1306 272414 20898
rect 271794 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 272414 -1306
rect 271794 -1626 272414 -1542
rect 271794 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 272414 -1626
rect 271794 -1894 272414 -1862
rect 275514 169174 276134 178000
rect 275514 168938 275546 169174
rect 275782 168938 275866 169174
rect 276102 168938 276134 169174
rect 275514 168854 276134 168938
rect 275514 168618 275546 168854
rect 275782 168618 275866 168854
rect 276102 168618 276134 168854
rect 275514 133174 276134 168618
rect 275514 132938 275546 133174
rect 275782 132938 275866 133174
rect 276102 132938 276134 133174
rect 275514 132854 276134 132938
rect 275514 132618 275546 132854
rect 275782 132618 275866 132854
rect 276102 132618 276134 132854
rect 275514 97174 276134 132618
rect 275514 96938 275546 97174
rect 275782 96938 275866 97174
rect 276102 96938 276134 97174
rect 275514 96854 276134 96938
rect 275514 96618 275546 96854
rect 275782 96618 275866 96854
rect 276102 96618 276134 96854
rect 275514 61174 276134 96618
rect 275514 60938 275546 61174
rect 275782 60938 275866 61174
rect 276102 60938 276134 61174
rect 275514 60854 276134 60938
rect 275514 60618 275546 60854
rect 275782 60618 275866 60854
rect 276102 60618 276134 60854
rect 275514 25174 276134 60618
rect 275514 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 276134 25174
rect 275514 24854 276134 24938
rect 275514 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 276134 24854
rect 275514 -3226 276134 24618
rect 275514 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 276134 -3226
rect 275514 -3546 276134 -3462
rect 275514 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 276134 -3546
rect 275514 -3814 276134 -3782
rect 279234 172894 279854 178000
rect 279234 172658 279266 172894
rect 279502 172658 279586 172894
rect 279822 172658 279854 172894
rect 279234 172574 279854 172658
rect 279234 172338 279266 172574
rect 279502 172338 279586 172574
rect 279822 172338 279854 172574
rect 279234 136894 279854 172338
rect 279234 136658 279266 136894
rect 279502 136658 279586 136894
rect 279822 136658 279854 136894
rect 279234 136574 279854 136658
rect 279234 136338 279266 136574
rect 279502 136338 279586 136574
rect 279822 136338 279854 136574
rect 279234 100894 279854 136338
rect 279234 100658 279266 100894
rect 279502 100658 279586 100894
rect 279822 100658 279854 100894
rect 279234 100574 279854 100658
rect 279234 100338 279266 100574
rect 279502 100338 279586 100574
rect 279822 100338 279854 100574
rect 279234 64894 279854 100338
rect 279234 64658 279266 64894
rect 279502 64658 279586 64894
rect 279822 64658 279854 64894
rect 279234 64574 279854 64658
rect 279234 64338 279266 64574
rect 279502 64338 279586 64574
rect 279822 64338 279854 64574
rect 279234 28894 279854 64338
rect 279234 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 279854 28894
rect 279234 28574 279854 28658
rect 279234 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 279854 28574
rect 279234 -5146 279854 28338
rect 279234 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 279854 -5146
rect 279234 -5466 279854 -5382
rect 279234 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 279854 -5466
rect 279234 -5734 279854 -5702
rect 282954 176614 283574 178000
rect 282954 176378 282986 176614
rect 283222 176378 283306 176614
rect 283542 176378 283574 176614
rect 282954 176294 283574 176378
rect 282954 176058 282986 176294
rect 283222 176058 283306 176294
rect 283542 176058 283574 176294
rect 282954 140614 283574 176058
rect 282954 140378 282986 140614
rect 283222 140378 283306 140614
rect 283542 140378 283574 140614
rect 282954 140294 283574 140378
rect 282954 140058 282986 140294
rect 283222 140058 283306 140294
rect 283542 140058 283574 140294
rect 282954 104614 283574 140058
rect 282954 104378 282986 104614
rect 283222 104378 283306 104614
rect 283542 104378 283574 104614
rect 282954 104294 283574 104378
rect 282954 104058 282986 104294
rect 283222 104058 283306 104294
rect 283542 104058 283574 104294
rect 282954 68614 283574 104058
rect 282954 68378 282986 68614
rect 283222 68378 283306 68614
rect 283542 68378 283574 68614
rect 282954 68294 283574 68378
rect 282954 68058 282986 68294
rect 283222 68058 283306 68294
rect 283542 68058 283574 68294
rect 282954 32614 283574 68058
rect 282954 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 283574 32614
rect 282954 32294 283574 32378
rect 282954 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 283574 32294
rect 264954 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 265574 -6106
rect 264954 -6426 265574 -6342
rect 264954 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 265574 -6426
rect 264954 -7654 265574 -6662
rect 282954 -7066 283574 32058
rect 289794 147454 290414 178000
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 289794 111454 290414 146898
rect 289794 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 290414 111454
rect 289794 111134 290414 111218
rect 289794 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 290414 111134
rect 289794 75454 290414 110898
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -1894 290414 -902
rect 293514 151174 294134 178000
rect 293514 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 294134 151174
rect 293514 150854 294134 150938
rect 293514 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 294134 150854
rect 293514 115174 294134 150618
rect 293514 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 294134 115174
rect 293514 114854 294134 114938
rect 293514 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 294134 114854
rect 293514 79174 294134 114618
rect 293514 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 294134 79174
rect 293514 78854 294134 78938
rect 293514 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 294134 78854
rect 293514 43174 294134 78618
rect 293514 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 294134 43174
rect 293514 42854 294134 42938
rect 293514 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 294134 42854
rect 293514 7174 294134 42618
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 293514 -2266 294134 6618
rect 293514 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 294134 -2266
rect 293514 -2586 294134 -2502
rect 293514 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 294134 -2586
rect 293514 -3814 294134 -2822
rect 297234 154894 297854 178000
rect 297234 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 297854 154894
rect 297234 154574 297854 154658
rect 297234 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 297854 154574
rect 297234 118894 297854 154338
rect 297234 118658 297266 118894
rect 297502 118658 297586 118894
rect 297822 118658 297854 118894
rect 297234 118574 297854 118658
rect 297234 118338 297266 118574
rect 297502 118338 297586 118574
rect 297822 118338 297854 118574
rect 297234 82894 297854 118338
rect 297234 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 297854 82894
rect 297234 82574 297854 82658
rect 297234 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 297854 82574
rect 297234 46894 297854 82338
rect 297234 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 297854 46894
rect 297234 46574 297854 46658
rect 297234 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 297854 46574
rect 297234 10894 297854 46338
rect 297234 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 297854 10894
rect 297234 10574 297854 10658
rect 297234 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 297854 10574
rect 297234 -4186 297854 10338
rect 297234 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 297854 -4186
rect 297234 -4506 297854 -4422
rect 297234 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 297854 -4506
rect 297234 -5734 297854 -4742
rect 300954 158614 301574 178000
rect 300954 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 301574 158614
rect 300954 158294 301574 158378
rect 300954 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 301574 158294
rect 300954 122614 301574 158058
rect 300954 122378 300986 122614
rect 301222 122378 301306 122614
rect 301542 122378 301574 122614
rect 300954 122294 301574 122378
rect 300954 122058 300986 122294
rect 301222 122058 301306 122294
rect 301542 122058 301574 122294
rect 300954 86614 301574 122058
rect 300954 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 301574 86614
rect 300954 86294 301574 86378
rect 300954 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 301574 86294
rect 300954 50614 301574 86058
rect 300954 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 301574 50614
rect 300954 50294 301574 50378
rect 300954 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 301574 50294
rect 300954 14614 301574 50058
rect 300954 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 301574 14614
rect 300954 14294 301574 14378
rect 300954 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 301574 14294
rect 282954 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 283574 -7066
rect 282954 -7386 283574 -7302
rect 282954 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 283574 -7386
rect 282954 -7654 283574 -7622
rect 300954 -6106 301574 14058
rect 307794 165454 308414 178000
rect 307794 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 308414 165454
rect 307794 165134 308414 165218
rect 307794 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 308414 165134
rect 307794 129454 308414 164898
rect 307794 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 308414 129454
rect 307794 129134 308414 129218
rect 307794 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 308414 129134
rect 307794 93454 308414 128898
rect 307794 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 308414 93454
rect 307794 93134 308414 93218
rect 307794 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 308414 93134
rect 307794 57454 308414 92898
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -1306 308414 20898
rect 307794 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 308414 -1306
rect 307794 -1626 308414 -1542
rect 307794 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 308414 -1626
rect 307794 -1894 308414 -1862
rect 311514 169174 312134 178000
rect 311514 168938 311546 169174
rect 311782 168938 311866 169174
rect 312102 168938 312134 169174
rect 311514 168854 312134 168938
rect 311514 168618 311546 168854
rect 311782 168618 311866 168854
rect 312102 168618 312134 168854
rect 311514 133174 312134 168618
rect 311514 132938 311546 133174
rect 311782 132938 311866 133174
rect 312102 132938 312134 133174
rect 311514 132854 312134 132938
rect 311514 132618 311546 132854
rect 311782 132618 311866 132854
rect 312102 132618 312134 132854
rect 311514 97174 312134 132618
rect 311514 96938 311546 97174
rect 311782 96938 311866 97174
rect 312102 96938 312134 97174
rect 311514 96854 312134 96938
rect 311514 96618 311546 96854
rect 311782 96618 311866 96854
rect 312102 96618 312134 96854
rect 311514 61174 312134 96618
rect 311514 60938 311546 61174
rect 311782 60938 311866 61174
rect 312102 60938 312134 61174
rect 311514 60854 312134 60938
rect 311514 60618 311546 60854
rect 311782 60618 311866 60854
rect 312102 60618 312134 60854
rect 311514 25174 312134 60618
rect 311514 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 312134 25174
rect 311514 24854 312134 24938
rect 311514 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 312134 24854
rect 311514 -3226 312134 24618
rect 311514 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 312134 -3226
rect 311514 -3546 312134 -3462
rect 311514 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 312134 -3546
rect 311514 -3814 312134 -3782
rect 315234 172894 315854 178000
rect 315234 172658 315266 172894
rect 315502 172658 315586 172894
rect 315822 172658 315854 172894
rect 315234 172574 315854 172658
rect 315234 172338 315266 172574
rect 315502 172338 315586 172574
rect 315822 172338 315854 172574
rect 315234 136894 315854 172338
rect 315234 136658 315266 136894
rect 315502 136658 315586 136894
rect 315822 136658 315854 136894
rect 315234 136574 315854 136658
rect 315234 136338 315266 136574
rect 315502 136338 315586 136574
rect 315822 136338 315854 136574
rect 315234 100894 315854 136338
rect 315234 100658 315266 100894
rect 315502 100658 315586 100894
rect 315822 100658 315854 100894
rect 315234 100574 315854 100658
rect 315234 100338 315266 100574
rect 315502 100338 315586 100574
rect 315822 100338 315854 100574
rect 315234 64894 315854 100338
rect 315234 64658 315266 64894
rect 315502 64658 315586 64894
rect 315822 64658 315854 64894
rect 315234 64574 315854 64658
rect 315234 64338 315266 64574
rect 315502 64338 315586 64574
rect 315822 64338 315854 64574
rect 315234 28894 315854 64338
rect 315234 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 315854 28894
rect 315234 28574 315854 28658
rect 315234 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 315854 28574
rect 315234 -5146 315854 28338
rect 315234 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 315854 -5146
rect 315234 -5466 315854 -5382
rect 315234 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 315854 -5466
rect 315234 -5734 315854 -5702
rect 318954 176614 319574 178000
rect 318954 176378 318986 176614
rect 319222 176378 319306 176614
rect 319542 176378 319574 176614
rect 318954 176294 319574 176378
rect 318954 176058 318986 176294
rect 319222 176058 319306 176294
rect 319542 176058 319574 176294
rect 318954 140614 319574 176058
rect 318954 140378 318986 140614
rect 319222 140378 319306 140614
rect 319542 140378 319574 140614
rect 318954 140294 319574 140378
rect 318954 140058 318986 140294
rect 319222 140058 319306 140294
rect 319542 140058 319574 140294
rect 318954 104614 319574 140058
rect 318954 104378 318986 104614
rect 319222 104378 319306 104614
rect 319542 104378 319574 104614
rect 318954 104294 319574 104378
rect 318954 104058 318986 104294
rect 319222 104058 319306 104294
rect 319542 104058 319574 104294
rect 318954 68614 319574 104058
rect 318954 68378 318986 68614
rect 319222 68378 319306 68614
rect 319542 68378 319574 68614
rect 318954 68294 319574 68378
rect 318954 68058 318986 68294
rect 319222 68058 319306 68294
rect 319542 68058 319574 68294
rect 318954 32614 319574 68058
rect 318954 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 319574 32614
rect 318954 32294 319574 32378
rect 318954 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 319574 32294
rect 300954 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 301574 -6106
rect 300954 -6426 301574 -6342
rect 300954 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 301574 -6426
rect 300954 -7654 301574 -6662
rect 318954 -7066 319574 32058
rect 325794 147454 326414 178000
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 325794 111454 326414 146898
rect 325794 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 326414 111454
rect 325794 111134 326414 111218
rect 325794 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 326414 111134
rect 325794 75454 326414 110898
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -1894 326414 -902
rect 329514 151174 330134 178000
rect 329514 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 330134 151174
rect 329514 150854 330134 150938
rect 329514 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 330134 150854
rect 329514 115174 330134 150618
rect 329514 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 330134 115174
rect 329514 114854 330134 114938
rect 329514 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 330134 114854
rect 329514 79174 330134 114618
rect 329514 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 330134 79174
rect 329514 78854 330134 78938
rect 329514 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 330134 78854
rect 329514 43174 330134 78618
rect 329514 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 330134 43174
rect 329514 42854 330134 42938
rect 329514 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 330134 42854
rect 329514 7174 330134 42618
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -2266 330134 6618
rect 329514 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 330134 -2266
rect 329514 -2586 330134 -2502
rect 329514 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 330134 -2586
rect 329514 -3814 330134 -2822
rect 333234 154894 333854 178000
rect 333234 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 333854 154894
rect 333234 154574 333854 154658
rect 333234 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 333854 154574
rect 333234 118894 333854 154338
rect 333234 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 333854 118894
rect 333234 118574 333854 118658
rect 333234 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 333854 118574
rect 333234 82894 333854 118338
rect 333234 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 333854 82894
rect 333234 82574 333854 82658
rect 333234 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 333854 82574
rect 333234 46894 333854 82338
rect 333234 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 333854 46894
rect 333234 46574 333854 46658
rect 333234 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 333854 46574
rect 333234 10894 333854 46338
rect 333234 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 333854 10894
rect 333234 10574 333854 10658
rect 333234 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 333854 10574
rect 333234 -4186 333854 10338
rect 333234 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 333854 -4186
rect 333234 -4506 333854 -4422
rect 333234 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 333854 -4506
rect 333234 -5734 333854 -4742
rect 336954 158614 337574 178000
rect 336954 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 337574 158614
rect 336954 158294 337574 158378
rect 336954 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 337574 158294
rect 336954 122614 337574 158058
rect 336954 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 337574 122614
rect 336954 122294 337574 122378
rect 336954 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 337574 122294
rect 336954 86614 337574 122058
rect 336954 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 337574 86614
rect 336954 86294 337574 86378
rect 336954 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 337574 86294
rect 336954 50614 337574 86058
rect 336954 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 337574 50614
rect 336954 50294 337574 50378
rect 336954 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 337574 50294
rect 336954 14614 337574 50058
rect 336954 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 337574 14614
rect 336954 14294 337574 14378
rect 336954 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 337574 14294
rect 318954 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 319574 -7066
rect 318954 -7386 319574 -7302
rect 318954 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 319574 -7386
rect 318954 -7654 319574 -7622
rect 336954 -6106 337574 14058
rect 343794 165454 344414 178000
rect 343794 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 344414 165454
rect 343794 165134 344414 165218
rect 343794 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 344414 165134
rect 343794 129454 344414 164898
rect 343794 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 344414 129454
rect 343794 129134 344414 129218
rect 343794 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 344414 129134
rect 343794 93454 344414 128898
rect 343794 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 344414 93454
rect 343794 93134 344414 93218
rect 343794 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 344414 93134
rect 343794 57454 344414 92898
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -1306 344414 20898
rect 343794 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 344414 -1306
rect 343794 -1626 344414 -1542
rect 343794 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 344414 -1626
rect 343794 -1894 344414 -1862
rect 347514 169174 348134 178000
rect 347514 168938 347546 169174
rect 347782 168938 347866 169174
rect 348102 168938 348134 169174
rect 347514 168854 348134 168938
rect 347514 168618 347546 168854
rect 347782 168618 347866 168854
rect 348102 168618 348134 168854
rect 347514 133174 348134 168618
rect 347514 132938 347546 133174
rect 347782 132938 347866 133174
rect 348102 132938 348134 133174
rect 347514 132854 348134 132938
rect 347514 132618 347546 132854
rect 347782 132618 347866 132854
rect 348102 132618 348134 132854
rect 347514 97174 348134 132618
rect 347514 96938 347546 97174
rect 347782 96938 347866 97174
rect 348102 96938 348134 97174
rect 347514 96854 348134 96938
rect 347514 96618 347546 96854
rect 347782 96618 347866 96854
rect 348102 96618 348134 96854
rect 347514 61174 348134 96618
rect 347514 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 348134 61174
rect 347514 60854 348134 60938
rect 347514 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 348134 60854
rect 347514 25174 348134 60618
rect 347514 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 348134 25174
rect 347514 24854 348134 24938
rect 347514 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 348134 24854
rect 347514 -3226 348134 24618
rect 347514 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 348134 -3226
rect 347514 -3546 348134 -3462
rect 347514 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 348134 -3546
rect 347514 -3814 348134 -3782
rect 351234 172894 351854 178000
rect 351234 172658 351266 172894
rect 351502 172658 351586 172894
rect 351822 172658 351854 172894
rect 351234 172574 351854 172658
rect 351234 172338 351266 172574
rect 351502 172338 351586 172574
rect 351822 172338 351854 172574
rect 351234 136894 351854 172338
rect 351234 136658 351266 136894
rect 351502 136658 351586 136894
rect 351822 136658 351854 136894
rect 351234 136574 351854 136658
rect 351234 136338 351266 136574
rect 351502 136338 351586 136574
rect 351822 136338 351854 136574
rect 351234 100894 351854 136338
rect 351234 100658 351266 100894
rect 351502 100658 351586 100894
rect 351822 100658 351854 100894
rect 351234 100574 351854 100658
rect 351234 100338 351266 100574
rect 351502 100338 351586 100574
rect 351822 100338 351854 100574
rect 351234 64894 351854 100338
rect 351234 64658 351266 64894
rect 351502 64658 351586 64894
rect 351822 64658 351854 64894
rect 351234 64574 351854 64658
rect 351234 64338 351266 64574
rect 351502 64338 351586 64574
rect 351822 64338 351854 64574
rect 351234 28894 351854 64338
rect 351234 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 351854 28894
rect 351234 28574 351854 28658
rect 351234 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 351854 28574
rect 351234 -5146 351854 28338
rect 351234 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 351854 -5146
rect 351234 -5466 351854 -5382
rect 351234 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 351854 -5466
rect 351234 -5734 351854 -5702
rect 354954 176614 355574 178000
rect 354954 176378 354986 176614
rect 355222 176378 355306 176614
rect 355542 176378 355574 176614
rect 354954 176294 355574 176378
rect 354954 176058 354986 176294
rect 355222 176058 355306 176294
rect 355542 176058 355574 176294
rect 354954 140614 355574 176058
rect 354954 140378 354986 140614
rect 355222 140378 355306 140614
rect 355542 140378 355574 140614
rect 354954 140294 355574 140378
rect 354954 140058 354986 140294
rect 355222 140058 355306 140294
rect 355542 140058 355574 140294
rect 354954 104614 355574 140058
rect 354954 104378 354986 104614
rect 355222 104378 355306 104614
rect 355542 104378 355574 104614
rect 354954 104294 355574 104378
rect 354954 104058 354986 104294
rect 355222 104058 355306 104294
rect 355542 104058 355574 104294
rect 354954 68614 355574 104058
rect 354954 68378 354986 68614
rect 355222 68378 355306 68614
rect 355542 68378 355574 68614
rect 354954 68294 355574 68378
rect 354954 68058 354986 68294
rect 355222 68058 355306 68294
rect 355542 68058 355574 68294
rect 354954 32614 355574 68058
rect 354954 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 355574 32614
rect 354954 32294 355574 32378
rect 354954 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 355574 32294
rect 336954 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 337574 -6106
rect 336954 -6426 337574 -6342
rect 336954 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 337574 -6426
rect 336954 -7654 337574 -6662
rect 354954 -7066 355574 32058
rect 361794 147454 362414 178000
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -1894 362414 -902
rect 365514 151174 366134 178000
rect 365514 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 366134 151174
rect 365514 150854 366134 150938
rect 365514 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 366134 150854
rect 365514 115174 366134 150618
rect 365514 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 366134 115174
rect 365514 114854 366134 114938
rect 365514 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 366134 114854
rect 365514 79174 366134 114618
rect 365514 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 366134 79174
rect 365514 78854 366134 78938
rect 365514 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 366134 78854
rect 365514 43174 366134 78618
rect 365514 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 366134 43174
rect 365514 42854 366134 42938
rect 365514 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 366134 42854
rect 365514 7174 366134 42618
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 365514 -2266 366134 6618
rect 365514 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 366134 -2266
rect 365514 -2586 366134 -2502
rect 365514 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 366134 -2586
rect 365514 -3814 366134 -2822
rect 369234 154894 369854 178000
rect 369234 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 369854 154894
rect 369234 154574 369854 154658
rect 369234 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 369854 154574
rect 369234 118894 369854 154338
rect 369234 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 369854 118894
rect 369234 118574 369854 118658
rect 369234 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 369854 118574
rect 369234 82894 369854 118338
rect 369234 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 369854 82894
rect 369234 82574 369854 82658
rect 369234 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 369854 82574
rect 369234 46894 369854 82338
rect 369234 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 369854 46894
rect 369234 46574 369854 46658
rect 369234 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 369854 46574
rect 369234 10894 369854 46338
rect 369234 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 369854 10894
rect 369234 10574 369854 10658
rect 369234 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 369854 10574
rect 369234 -4186 369854 10338
rect 369234 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 369854 -4186
rect 369234 -4506 369854 -4422
rect 369234 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 369854 -4506
rect 369234 -5734 369854 -4742
rect 372954 158614 373574 178000
rect 372954 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 373574 158614
rect 372954 158294 373574 158378
rect 372954 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 373574 158294
rect 372954 122614 373574 158058
rect 372954 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 373574 122614
rect 372954 122294 373574 122378
rect 372954 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 373574 122294
rect 372954 86614 373574 122058
rect 372954 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 373574 86614
rect 372954 86294 373574 86378
rect 372954 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 373574 86294
rect 372954 50614 373574 86058
rect 372954 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 373574 50614
rect 372954 50294 373574 50378
rect 372954 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 373574 50294
rect 372954 14614 373574 50058
rect 372954 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 373574 14614
rect 372954 14294 373574 14378
rect 372954 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 373574 14294
rect 354954 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 355574 -7066
rect 354954 -7386 355574 -7302
rect 354954 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 355574 -7386
rect 354954 -7654 355574 -7622
rect 372954 -6106 373574 14058
rect 379794 165454 380414 178000
rect 379794 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 380414 165454
rect 379794 165134 380414 165218
rect 379794 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 380414 165134
rect 379794 129454 380414 164898
rect 379794 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 380414 129454
rect 379794 129134 380414 129218
rect 379794 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 380414 129134
rect 379794 93454 380414 128898
rect 379794 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 380414 93454
rect 379794 93134 380414 93218
rect 379794 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 380414 93134
rect 379794 57454 380414 92898
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -1306 380414 20898
rect 379794 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 380414 -1306
rect 379794 -1626 380414 -1542
rect 379794 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 380414 -1626
rect 379794 -1894 380414 -1862
rect 383514 169174 384134 178000
rect 383514 168938 383546 169174
rect 383782 168938 383866 169174
rect 384102 168938 384134 169174
rect 383514 168854 384134 168938
rect 383514 168618 383546 168854
rect 383782 168618 383866 168854
rect 384102 168618 384134 168854
rect 383514 133174 384134 168618
rect 383514 132938 383546 133174
rect 383782 132938 383866 133174
rect 384102 132938 384134 133174
rect 383514 132854 384134 132938
rect 383514 132618 383546 132854
rect 383782 132618 383866 132854
rect 384102 132618 384134 132854
rect 383514 97174 384134 132618
rect 383514 96938 383546 97174
rect 383782 96938 383866 97174
rect 384102 96938 384134 97174
rect 383514 96854 384134 96938
rect 383514 96618 383546 96854
rect 383782 96618 383866 96854
rect 384102 96618 384134 96854
rect 383514 61174 384134 96618
rect 383514 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 384134 61174
rect 383514 60854 384134 60938
rect 383514 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 384134 60854
rect 383514 25174 384134 60618
rect 383514 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 384134 25174
rect 383514 24854 384134 24938
rect 383514 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 384134 24854
rect 383514 -3226 384134 24618
rect 383514 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 384134 -3226
rect 383514 -3546 384134 -3462
rect 383514 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 384134 -3546
rect 383514 -3814 384134 -3782
rect 387234 172894 387854 178000
rect 387234 172658 387266 172894
rect 387502 172658 387586 172894
rect 387822 172658 387854 172894
rect 387234 172574 387854 172658
rect 387234 172338 387266 172574
rect 387502 172338 387586 172574
rect 387822 172338 387854 172574
rect 387234 136894 387854 172338
rect 387234 136658 387266 136894
rect 387502 136658 387586 136894
rect 387822 136658 387854 136894
rect 387234 136574 387854 136658
rect 387234 136338 387266 136574
rect 387502 136338 387586 136574
rect 387822 136338 387854 136574
rect 387234 100894 387854 136338
rect 387234 100658 387266 100894
rect 387502 100658 387586 100894
rect 387822 100658 387854 100894
rect 387234 100574 387854 100658
rect 387234 100338 387266 100574
rect 387502 100338 387586 100574
rect 387822 100338 387854 100574
rect 387234 64894 387854 100338
rect 387234 64658 387266 64894
rect 387502 64658 387586 64894
rect 387822 64658 387854 64894
rect 387234 64574 387854 64658
rect 387234 64338 387266 64574
rect 387502 64338 387586 64574
rect 387822 64338 387854 64574
rect 387234 28894 387854 64338
rect 387234 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 387854 28894
rect 387234 28574 387854 28658
rect 387234 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 387854 28574
rect 387234 -5146 387854 28338
rect 387234 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 387854 -5146
rect 387234 -5466 387854 -5382
rect 387234 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 387854 -5466
rect 387234 -5734 387854 -5702
rect 390954 176614 391574 178000
rect 390954 176378 390986 176614
rect 391222 176378 391306 176614
rect 391542 176378 391574 176614
rect 390954 176294 391574 176378
rect 390954 176058 390986 176294
rect 391222 176058 391306 176294
rect 391542 176058 391574 176294
rect 390954 140614 391574 176058
rect 390954 140378 390986 140614
rect 391222 140378 391306 140614
rect 391542 140378 391574 140614
rect 390954 140294 391574 140378
rect 390954 140058 390986 140294
rect 391222 140058 391306 140294
rect 391542 140058 391574 140294
rect 390954 104614 391574 140058
rect 390954 104378 390986 104614
rect 391222 104378 391306 104614
rect 391542 104378 391574 104614
rect 390954 104294 391574 104378
rect 390954 104058 390986 104294
rect 391222 104058 391306 104294
rect 391542 104058 391574 104294
rect 390954 68614 391574 104058
rect 390954 68378 390986 68614
rect 391222 68378 391306 68614
rect 391542 68378 391574 68614
rect 390954 68294 391574 68378
rect 390954 68058 390986 68294
rect 391222 68058 391306 68294
rect 391542 68058 391574 68294
rect 390954 32614 391574 68058
rect 390954 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 391574 32614
rect 390954 32294 391574 32378
rect 390954 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 391574 32294
rect 372954 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 373574 -6106
rect 372954 -6426 373574 -6342
rect 372954 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 373574 -6426
rect 372954 -7654 373574 -6662
rect 390954 -7066 391574 32058
rect 397794 147454 398414 178000
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -1894 398414 -902
rect 401514 151174 402134 178000
rect 401514 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 402134 151174
rect 401514 150854 402134 150938
rect 401514 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 402134 150854
rect 401514 115174 402134 150618
rect 401514 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 402134 115174
rect 401514 114854 402134 114938
rect 401514 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 402134 114854
rect 401514 79174 402134 114618
rect 401514 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 402134 79174
rect 401514 78854 402134 78938
rect 401514 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 402134 78854
rect 401514 43174 402134 78618
rect 401514 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 402134 43174
rect 401514 42854 402134 42938
rect 401514 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 402134 42854
rect 401514 7174 402134 42618
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -2266 402134 6618
rect 401514 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 402134 -2266
rect 401514 -2586 402134 -2502
rect 401514 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 402134 -2586
rect 401514 -3814 402134 -2822
rect 405234 154894 405854 178000
rect 405234 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 405854 154894
rect 405234 154574 405854 154658
rect 405234 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 405854 154574
rect 405234 118894 405854 154338
rect 405234 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 405854 118894
rect 405234 118574 405854 118658
rect 405234 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 405854 118574
rect 405234 82894 405854 118338
rect 405234 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 405854 82894
rect 405234 82574 405854 82658
rect 405234 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 405854 82574
rect 405234 46894 405854 82338
rect 405234 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 405854 46894
rect 405234 46574 405854 46658
rect 405234 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 405854 46574
rect 405234 10894 405854 46338
rect 405234 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 405854 10894
rect 405234 10574 405854 10658
rect 405234 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 405854 10574
rect 405234 -4186 405854 10338
rect 405234 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 405854 -4186
rect 405234 -4506 405854 -4422
rect 405234 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 405854 -4506
rect 405234 -5734 405854 -4742
rect 408954 158614 409574 178000
rect 408954 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 409574 158614
rect 408954 158294 409574 158378
rect 408954 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 409574 158294
rect 408954 122614 409574 158058
rect 408954 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 409574 122614
rect 408954 122294 409574 122378
rect 408954 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 409574 122294
rect 408954 86614 409574 122058
rect 408954 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 409574 86614
rect 408954 86294 409574 86378
rect 408954 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 409574 86294
rect 408954 50614 409574 86058
rect 408954 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 409574 50614
rect 408954 50294 409574 50378
rect 408954 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 409574 50294
rect 408954 14614 409574 50058
rect 408954 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 409574 14614
rect 408954 14294 409574 14378
rect 408954 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 409574 14294
rect 390954 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 391574 -7066
rect 390954 -7386 391574 -7302
rect 390954 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 391574 -7386
rect 390954 -7654 391574 -7622
rect 408954 -6106 409574 14058
rect 415794 165454 416414 178000
rect 415794 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 416414 165454
rect 415794 165134 416414 165218
rect 415794 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 416414 165134
rect 415794 129454 416414 164898
rect 415794 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 416414 129454
rect 415794 129134 416414 129218
rect 415794 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 416414 129134
rect 415794 93454 416414 128898
rect 415794 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 416414 93454
rect 415794 93134 416414 93218
rect 415794 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 416414 93134
rect 415794 57454 416414 92898
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -1306 416414 20898
rect 415794 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 416414 -1306
rect 415794 -1626 416414 -1542
rect 415794 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 416414 -1626
rect 415794 -1894 416414 -1862
rect 419514 169174 420134 178000
rect 419514 168938 419546 169174
rect 419782 168938 419866 169174
rect 420102 168938 420134 169174
rect 419514 168854 420134 168938
rect 419514 168618 419546 168854
rect 419782 168618 419866 168854
rect 420102 168618 420134 168854
rect 419514 133174 420134 168618
rect 419514 132938 419546 133174
rect 419782 132938 419866 133174
rect 420102 132938 420134 133174
rect 419514 132854 420134 132938
rect 419514 132618 419546 132854
rect 419782 132618 419866 132854
rect 420102 132618 420134 132854
rect 419514 97174 420134 132618
rect 419514 96938 419546 97174
rect 419782 96938 419866 97174
rect 420102 96938 420134 97174
rect 419514 96854 420134 96938
rect 419514 96618 419546 96854
rect 419782 96618 419866 96854
rect 420102 96618 420134 96854
rect 419514 61174 420134 96618
rect 419514 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 420134 61174
rect 419514 60854 420134 60938
rect 419514 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 420134 60854
rect 419514 25174 420134 60618
rect 419514 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 420134 25174
rect 419514 24854 420134 24938
rect 419514 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 420134 24854
rect 419514 -3226 420134 24618
rect 419514 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 420134 -3226
rect 419514 -3546 420134 -3462
rect 419514 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 420134 -3546
rect 419514 -3814 420134 -3782
rect 423234 172894 423854 178000
rect 423234 172658 423266 172894
rect 423502 172658 423586 172894
rect 423822 172658 423854 172894
rect 423234 172574 423854 172658
rect 423234 172338 423266 172574
rect 423502 172338 423586 172574
rect 423822 172338 423854 172574
rect 423234 136894 423854 172338
rect 423234 136658 423266 136894
rect 423502 136658 423586 136894
rect 423822 136658 423854 136894
rect 423234 136574 423854 136658
rect 423234 136338 423266 136574
rect 423502 136338 423586 136574
rect 423822 136338 423854 136574
rect 423234 100894 423854 136338
rect 423234 100658 423266 100894
rect 423502 100658 423586 100894
rect 423822 100658 423854 100894
rect 423234 100574 423854 100658
rect 423234 100338 423266 100574
rect 423502 100338 423586 100574
rect 423822 100338 423854 100574
rect 423234 64894 423854 100338
rect 423234 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 423854 64894
rect 423234 64574 423854 64658
rect 423234 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 423854 64574
rect 423234 28894 423854 64338
rect 423234 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 423854 28894
rect 423234 28574 423854 28658
rect 423234 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 423854 28574
rect 423234 -5146 423854 28338
rect 423234 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 423854 -5146
rect 423234 -5466 423854 -5382
rect 423234 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 423854 -5466
rect 423234 -5734 423854 -5702
rect 426954 176614 427574 178000
rect 426954 176378 426986 176614
rect 427222 176378 427306 176614
rect 427542 176378 427574 176614
rect 426954 176294 427574 176378
rect 426954 176058 426986 176294
rect 427222 176058 427306 176294
rect 427542 176058 427574 176294
rect 426954 140614 427574 176058
rect 426954 140378 426986 140614
rect 427222 140378 427306 140614
rect 427542 140378 427574 140614
rect 426954 140294 427574 140378
rect 426954 140058 426986 140294
rect 427222 140058 427306 140294
rect 427542 140058 427574 140294
rect 426954 104614 427574 140058
rect 426954 104378 426986 104614
rect 427222 104378 427306 104614
rect 427542 104378 427574 104614
rect 426954 104294 427574 104378
rect 426954 104058 426986 104294
rect 427222 104058 427306 104294
rect 427542 104058 427574 104294
rect 426954 68614 427574 104058
rect 426954 68378 426986 68614
rect 427222 68378 427306 68614
rect 427542 68378 427574 68614
rect 426954 68294 427574 68378
rect 426954 68058 426986 68294
rect 427222 68058 427306 68294
rect 427542 68058 427574 68294
rect 426954 32614 427574 68058
rect 426954 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 427574 32614
rect 426954 32294 427574 32378
rect 426954 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 427574 32294
rect 408954 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 409574 -6106
rect 408954 -6426 409574 -6342
rect 408954 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 409574 -6426
rect 408954 -7654 409574 -6662
rect 426954 -7066 427574 32058
rect 433794 147454 434414 178000
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 111454 434414 146898
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -1894 434414 -902
rect 437514 151174 438134 178000
rect 437514 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 438134 151174
rect 437514 150854 438134 150938
rect 437514 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 438134 150854
rect 437514 115174 438134 150618
rect 437514 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 438134 115174
rect 437514 114854 438134 114938
rect 437514 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 438134 114854
rect 437514 79174 438134 114618
rect 437514 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 438134 79174
rect 437514 78854 438134 78938
rect 437514 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 438134 78854
rect 437514 43174 438134 78618
rect 437514 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 438134 43174
rect 437514 42854 438134 42938
rect 437514 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 438134 42854
rect 437514 7174 438134 42618
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -2266 438134 6618
rect 437514 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 438134 -2266
rect 437514 -2586 438134 -2502
rect 437514 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 438134 -2586
rect 437514 -3814 438134 -2822
rect 441234 154894 441854 178000
rect 441234 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 441854 154894
rect 441234 154574 441854 154658
rect 441234 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 441854 154574
rect 441234 118894 441854 154338
rect 441234 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 441854 118894
rect 441234 118574 441854 118658
rect 441234 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 441854 118574
rect 441234 82894 441854 118338
rect 441234 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 441854 82894
rect 441234 82574 441854 82658
rect 441234 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 441854 82574
rect 441234 46894 441854 82338
rect 441234 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 441854 46894
rect 441234 46574 441854 46658
rect 441234 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 441854 46574
rect 441234 10894 441854 46338
rect 441234 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 441854 10894
rect 441234 10574 441854 10658
rect 441234 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 441854 10574
rect 441234 -4186 441854 10338
rect 441234 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 441854 -4186
rect 441234 -4506 441854 -4422
rect 441234 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 441854 -4506
rect 441234 -5734 441854 -4742
rect 444954 158614 445574 178000
rect 444954 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 445574 158614
rect 444954 158294 445574 158378
rect 444954 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 445574 158294
rect 444954 122614 445574 158058
rect 444954 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 445574 122614
rect 444954 122294 445574 122378
rect 444954 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 445574 122294
rect 444954 86614 445574 122058
rect 444954 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 445574 86614
rect 444954 86294 445574 86378
rect 444954 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 445574 86294
rect 444954 50614 445574 86058
rect 444954 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 445574 50614
rect 444954 50294 445574 50378
rect 444954 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 445574 50294
rect 444954 14614 445574 50058
rect 444954 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 445574 14614
rect 444954 14294 445574 14378
rect 444954 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 445574 14294
rect 426954 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 427574 -7066
rect 426954 -7386 427574 -7302
rect 426954 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 427574 -7386
rect 426954 -7654 427574 -7622
rect 444954 -6106 445574 14058
rect 451794 165454 452414 178000
rect 451794 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 452414 165454
rect 451794 165134 452414 165218
rect 451794 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 452414 165134
rect 451794 129454 452414 164898
rect 451794 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 452414 129454
rect 451794 129134 452414 129218
rect 451794 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 452414 129134
rect 451794 93454 452414 128898
rect 451794 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 452414 93454
rect 451794 93134 452414 93218
rect 451794 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 452414 93134
rect 451794 57454 452414 92898
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -1306 452414 20898
rect 451794 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 452414 -1306
rect 451794 -1626 452414 -1542
rect 451794 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 452414 -1626
rect 451794 -1894 452414 -1862
rect 455514 169174 456134 178000
rect 455514 168938 455546 169174
rect 455782 168938 455866 169174
rect 456102 168938 456134 169174
rect 455514 168854 456134 168938
rect 455514 168618 455546 168854
rect 455782 168618 455866 168854
rect 456102 168618 456134 168854
rect 455514 133174 456134 168618
rect 455514 132938 455546 133174
rect 455782 132938 455866 133174
rect 456102 132938 456134 133174
rect 455514 132854 456134 132938
rect 455514 132618 455546 132854
rect 455782 132618 455866 132854
rect 456102 132618 456134 132854
rect 455514 97174 456134 132618
rect 455514 96938 455546 97174
rect 455782 96938 455866 97174
rect 456102 96938 456134 97174
rect 455514 96854 456134 96938
rect 455514 96618 455546 96854
rect 455782 96618 455866 96854
rect 456102 96618 456134 96854
rect 455514 61174 456134 96618
rect 455514 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 456134 61174
rect 455514 60854 456134 60938
rect 455514 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 456134 60854
rect 455514 25174 456134 60618
rect 455514 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 456134 25174
rect 455514 24854 456134 24938
rect 455514 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 456134 24854
rect 455514 -3226 456134 24618
rect 455514 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 456134 -3226
rect 455514 -3546 456134 -3462
rect 455514 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 456134 -3546
rect 455514 -3814 456134 -3782
rect 459234 172894 459854 178000
rect 459234 172658 459266 172894
rect 459502 172658 459586 172894
rect 459822 172658 459854 172894
rect 459234 172574 459854 172658
rect 459234 172338 459266 172574
rect 459502 172338 459586 172574
rect 459822 172338 459854 172574
rect 459234 136894 459854 172338
rect 459234 136658 459266 136894
rect 459502 136658 459586 136894
rect 459822 136658 459854 136894
rect 459234 136574 459854 136658
rect 459234 136338 459266 136574
rect 459502 136338 459586 136574
rect 459822 136338 459854 136574
rect 459234 100894 459854 136338
rect 459234 100658 459266 100894
rect 459502 100658 459586 100894
rect 459822 100658 459854 100894
rect 459234 100574 459854 100658
rect 459234 100338 459266 100574
rect 459502 100338 459586 100574
rect 459822 100338 459854 100574
rect 459234 64894 459854 100338
rect 459234 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 459854 64894
rect 459234 64574 459854 64658
rect 459234 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 459854 64574
rect 459234 28894 459854 64338
rect 459234 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 459854 28894
rect 459234 28574 459854 28658
rect 459234 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 459854 28574
rect 459234 -5146 459854 28338
rect 459234 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 459854 -5146
rect 459234 -5466 459854 -5382
rect 459234 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 459854 -5466
rect 459234 -5734 459854 -5702
rect 462954 176614 463574 178000
rect 462954 176378 462986 176614
rect 463222 176378 463306 176614
rect 463542 176378 463574 176614
rect 462954 176294 463574 176378
rect 462954 176058 462986 176294
rect 463222 176058 463306 176294
rect 463542 176058 463574 176294
rect 462954 140614 463574 176058
rect 462954 140378 462986 140614
rect 463222 140378 463306 140614
rect 463542 140378 463574 140614
rect 462954 140294 463574 140378
rect 462954 140058 462986 140294
rect 463222 140058 463306 140294
rect 463542 140058 463574 140294
rect 462954 104614 463574 140058
rect 462954 104378 462986 104614
rect 463222 104378 463306 104614
rect 463542 104378 463574 104614
rect 462954 104294 463574 104378
rect 462954 104058 462986 104294
rect 463222 104058 463306 104294
rect 463542 104058 463574 104294
rect 462954 68614 463574 104058
rect 462954 68378 462986 68614
rect 463222 68378 463306 68614
rect 463542 68378 463574 68614
rect 462954 68294 463574 68378
rect 462954 68058 462986 68294
rect 463222 68058 463306 68294
rect 463542 68058 463574 68294
rect 462954 32614 463574 68058
rect 462954 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 463574 32614
rect 462954 32294 463574 32378
rect 462954 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 463574 32294
rect 444954 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 445574 -6106
rect 444954 -6426 445574 -6342
rect 444954 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 445574 -6426
rect 444954 -7654 445574 -6662
rect 462954 -7066 463574 32058
rect 469794 147454 470414 178000
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -1894 470414 -902
rect 473514 151174 474134 178000
rect 473514 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 474134 151174
rect 473514 150854 474134 150938
rect 473514 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 474134 150854
rect 473514 115174 474134 150618
rect 473514 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 474134 115174
rect 473514 114854 474134 114938
rect 473514 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 474134 114854
rect 473514 79174 474134 114618
rect 473514 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 474134 79174
rect 473514 78854 474134 78938
rect 473514 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 474134 78854
rect 473514 43174 474134 78618
rect 473514 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 474134 43174
rect 473514 42854 474134 42938
rect 473514 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 474134 42854
rect 473514 7174 474134 42618
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -2266 474134 6618
rect 473514 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 474134 -2266
rect 473514 -2586 474134 -2502
rect 473514 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 474134 -2586
rect 473514 -3814 474134 -2822
rect 477234 154894 477854 178000
rect 477234 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 477854 154894
rect 477234 154574 477854 154658
rect 477234 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 477854 154574
rect 477234 118894 477854 154338
rect 477234 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 477854 118894
rect 477234 118574 477854 118658
rect 477234 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 477854 118574
rect 477234 82894 477854 118338
rect 477234 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 477854 82894
rect 477234 82574 477854 82658
rect 477234 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 477854 82574
rect 477234 46894 477854 82338
rect 477234 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 477854 46894
rect 477234 46574 477854 46658
rect 477234 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 477854 46574
rect 477234 10894 477854 46338
rect 477234 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 477854 10894
rect 477234 10574 477854 10658
rect 477234 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 477854 10574
rect 477234 -4186 477854 10338
rect 477234 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 477854 -4186
rect 477234 -4506 477854 -4422
rect 477234 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 477854 -4506
rect 477234 -5734 477854 -4742
rect 480954 158614 481574 178000
rect 480954 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 481574 158614
rect 480954 158294 481574 158378
rect 480954 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 481574 158294
rect 480954 122614 481574 158058
rect 480954 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 481574 122614
rect 480954 122294 481574 122378
rect 480954 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 481574 122294
rect 480954 86614 481574 122058
rect 480954 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 481574 86614
rect 480954 86294 481574 86378
rect 480954 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 481574 86294
rect 480954 50614 481574 86058
rect 480954 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 481574 50614
rect 480954 50294 481574 50378
rect 480954 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 481574 50294
rect 480954 14614 481574 50058
rect 480954 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 481574 14614
rect 480954 14294 481574 14378
rect 480954 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 481574 14294
rect 462954 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 463574 -7066
rect 462954 -7386 463574 -7302
rect 462954 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 463574 -7386
rect 462954 -7654 463574 -7622
rect 480954 -6106 481574 14058
rect 487794 165454 488414 178000
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 129454 488414 164898
rect 487794 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 488414 129454
rect 487794 129134 488414 129218
rect 487794 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 488414 129134
rect 487794 93454 488414 128898
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -1306 488414 20898
rect 487794 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 488414 -1306
rect 487794 -1626 488414 -1542
rect 487794 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 488414 -1626
rect 487794 -1894 488414 -1862
rect 491514 169174 492134 178000
rect 491514 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 492134 169174
rect 491514 168854 492134 168938
rect 491514 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 492134 168854
rect 491514 133174 492134 168618
rect 491514 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 492134 133174
rect 491514 132854 492134 132938
rect 491514 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 492134 132854
rect 491514 97174 492134 132618
rect 491514 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 492134 97174
rect 491514 96854 492134 96938
rect 491514 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 492134 96854
rect 491514 61174 492134 96618
rect 491514 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 492134 61174
rect 491514 60854 492134 60938
rect 491514 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 492134 60854
rect 491514 25174 492134 60618
rect 491514 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 492134 25174
rect 491514 24854 492134 24938
rect 491514 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 492134 24854
rect 491514 -3226 492134 24618
rect 491514 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 492134 -3226
rect 491514 -3546 492134 -3462
rect 491514 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 492134 -3546
rect 491514 -3814 492134 -3782
rect 495234 172894 495854 178000
rect 495234 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 495854 172894
rect 495234 172574 495854 172658
rect 495234 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 495854 172574
rect 495234 136894 495854 172338
rect 495234 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 495854 136894
rect 495234 136574 495854 136658
rect 495234 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 495854 136574
rect 495234 100894 495854 136338
rect 495234 100658 495266 100894
rect 495502 100658 495586 100894
rect 495822 100658 495854 100894
rect 495234 100574 495854 100658
rect 495234 100338 495266 100574
rect 495502 100338 495586 100574
rect 495822 100338 495854 100574
rect 495234 64894 495854 100338
rect 495234 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 495854 64894
rect 495234 64574 495854 64658
rect 495234 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 495854 64574
rect 495234 28894 495854 64338
rect 495234 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 495854 28894
rect 495234 28574 495854 28658
rect 495234 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 495854 28574
rect 495234 -5146 495854 28338
rect 495234 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 495854 -5146
rect 495234 -5466 495854 -5382
rect 495234 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 495854 -5466
rect 495234 -5734 495854 -5702
rect 498954 176614 499574 178000
rect 498954 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 499574 176614
rect 498954 176294 499574 176378
rect 498954 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 499574 176294
rect 498954 140614 499574 176058
rect 498954 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 499574 140614
rect 498954 140294 499574 140378
rect 498954 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 499574 140294
rect 498954 104614 499574 140058
rect 498954 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 499574 104614
rect 498954 104294 499574 104378
rect 498954 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 499574 104294
rect 498954 68614 499574 104058
rect 498954 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 499574 68614
rect 498954 68294 499574 68378
rect 498954 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 499574 68294
rect 498954 32614 499574 68058
rect 498954 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 499574 32614
rect 498954 32294 499574 32378
rect 498954 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 499574 32294
rect 480954 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 481574 -6106
rect 480954 -6426 481574 -6342
rect 480954 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 481574 -6426
rect 480954 -7654 481574 -6662
rect 498954 -7066 499574 32058
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -1894 506414 -902
rect 509514 691174 510134 706202
rect 509514 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 510134 691174
rect 509514 690854 510134 690938
rect 509514 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 510134 690854
rect 509514 655174 510134 690618
rect 509514 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 510134 655174
rect 509514 654854 510134 654938
rect 509514 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 510134 654854
rect 509514 619174 510134 654618
rect 509514 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 510134 619174
rect 509514 618854 510134 618938
rect 509514 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 510134 618854
rect 509514 583174 510134 618618
rect 509514 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 510134 583174
rect 509514 582854 510134 582938
rect 509514 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 510134 582854
rect 509514 547174 510134 582618
rect 509514 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 510134 547174
rect 509514 546854 510134 546938
rect 509514 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 510134 546854
rect 509514 511174 510134 546618
rect 509514 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 510134 511174
rect 509514 510854 510134 510938
rect 509514 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 510134 510854
rect 509514 475174 510134 510618
rect 509514 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 510134 475174
rect 509514 474854 510134 474938
rect 509514 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 510134 474854
rect 509514 439174 510134 474618
rect 509514 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 510134 439174
rect 509514 438854 510134 438938
rect 509514 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 510134 438854
rect 509514 403174 510134 438618
rect 509514 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 510134 403174
rect 509514 402854 510134 402938
rect 509514 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 510134 402854
rect 509514 367174 510134 402618
rect 509514 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 510134 367174
rect 509514 366854 510134 366938
rect 509514 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 510134 366854
rect 509514 331174 510134 366618
rect 509514 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 510134 331174
rect 509514 330854 510134 330938
rect 509514 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 510134 330854
rect 509514 295174 510134 330618
rect 509514 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 510134 295174
rect 509514 294854 510134 294938
rect 509514 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 510134 294854
rect 509514 259174 510134 294618
rect 509514 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 510134 259174
rect 509514 258854 510134 258938
rect 509514 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 510134 258854
rect 509514 223174 510134 258618
rect 509514 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 510134 223174
rect 509514 222854 510134 222938
rect 509514 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 510134 222854
rect 509514 187174 510134 222618
rect 509514 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 510134 187174
rect 509514 186854 510134 186938
rect 509514 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 510134 186854
rect 509514 151174 510134 186618
rect 509514 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 510134 151174
rect 509514 150854 510134 150938
rect 509514 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 510134 150854
rect 509514 115174 510134 150618
rect 509514 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 510134 115174
rect 509514 114854 510134 114938
rect 509514 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 510134 114854
rect 509514 79174 510134 114618
rect 509514 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 510134 79174
rect 509514 78854 510134 78938
rect 509514 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 510134 78854
rect 509514 43174 510134 78618
rect 509514 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 510134 43174
rect 509514 42854 510134 42938
rect 509514 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 510134 42854
rect 509514 7174 510134 42618
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -2266 510134 6618
rect 509514 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 510134 -2266
rect 509514 -2586 510134 -2502
rect 509514 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 510134 -2586
rect 509514 -3814 510134 -2822
rect 513234 694894 513854 708122
rect 513234 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 513854 694894
rect 513234 694574 513854 694658
rect 513234 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 513854 694574
rect 513234 658894 513854 694338
rect 513234 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 513854 658894
rect 513234 658574 513854 658658
rect 513234 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 513854 658574
rect 513234 622894 513854 658338
rect 513234 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 513854 622894
rect 513234 622574 513854 622658
rect 513234 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 513854 622574
rect 513234 586894 513854 622338
rect 513234 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 513854 586894
rect 513234 586574 513854 586658
rect 513234 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 513854 586574
rect 513234 550894 513854 586338
rect 513234 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 513854 550894
rect 513234 550574 513854 550658
rect 513234 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 513854 550574
rect 513234 514894 513854 550338
rect 513234 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 513854 514894
rect 513234 514574 513854 514658
rect 513234 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 513854 514574
rect 513234 478894 513854 514338
rect 513234 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 513854 478894
rect 513234 478574 513854 478658
rect 513234 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 513854 478574
rect 513234 442894 513854 478338
rect 513234 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 513854 442894
rect 513234 442574 513854 442658
rect 513234 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 513854 442574
rect 513234 406894 513854 442338
rect 513234 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 513854 406894
rect 513234 406574 513854 406658
rect 513234 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 513854 406574
rect 513234 370894 513854 406338
rect 513234 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 513854 370894
rect 513234 370574 513854 370658
rect 513234 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 513854 370574
rect 513234 334894 513854 370338
rect 513234 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 513854 334894
rect 513234 334574 513854 334658
rect 513234 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 513854 334574
rect 513234 298894 513854 334338
rect 513234 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 513854 298894
rect 513234 298574 513854 298658
rect 513234 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 513854 298574
rect 513234 262894 513854 298338
rect 513234 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 513854 262894
rect 513234 262574 513854 262658
rect 513234 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 513854 262574
rect 513234 226894 513854 262338
rect 513234 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 513854 226894
rect 513234 226574 513854 226658
rect 513234 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 513854 226574
rect 513234 190894 513854 226338
rect 513234 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 513854 190894
rect 513234 190574 513854 190658
rect 513234 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 513854 190574
rect 513234 154894 513854 190338
rect 513234 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 513854 154894
rect 513234 154574 513854 154658
rect 513234 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 513854 154574
rect 513234 118894 513854 154338
rect 513234 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 513854 118894
rect 513234 118574 513854 118658
rect 513234 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 513854 118574
rect 513234 82894 513854 118338
rect 513234 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 513854 82894
rect 513234 82574 513854 82658
rect 513234 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 513854 82574
rect 513234 46894 513854 82338
rect 513234 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 513854 46894
rect 513234 46574 513854 46658
rect 513234 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 513854 46574
rect 513234 10894 513854 46338
rect 513234 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 513854 10894
rect 513234 10574 513854 10658
rect 513234 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 513854 10574
rect 513234 -4186 513854 10338
rect 513234 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 513854 -4186
rect 513234 -4506 513854 -4422
rect 513234 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 513854 -4506
rect 513234 -5734 513854 -4742
rect 516954 698614 517574 710042
rect 534954 711558 535574 711590
rect 534954 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 535574 711558
rect 534954 711238 535574 711322
rect 534954 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 535574 711238
rect 531234 709638 531854 709670
rect 531234 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 531854 709638
rect 531234 709318 531854 709402
rect 531234 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 531854 709318
rect 527514 707718 528134 707750
rect 527514 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 528134 707718
rect 527514 707398 528134 707482
rect 527514 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 528134 707398
rect 516954 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 517574 698614
rect 516954 698294 517574 698378
rect 516954 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 517574 698294
rect 516954 662614 517574 698058
rect 516954 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 517574 662614
rect 516954 662294 517574 662378
rect 516954 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 517574 662294
rect 516954 626614 517574 662058
rect 516954 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 517574 626614
rect 516954 626294 517574 626378
rect 516954 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 517574 626294
rect 516954 590614 517574 626058
rect 516954 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 517574 590614
rect 516954 590294 517574 590378
rect 516954 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 517574 590294
rect 516954 554614 517574 590058
rect 516954 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 517574 554614
rect 516954 554294 517574 554378
rect 516954 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 517574 554294
rect 516954 518614 517574 554058
rect 516954 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 517574 518614
rect 516954 518294 517574 518378
rect 516954 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 517574 518294
rect 516954 482614 517574 518058
rect 516954 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 517574 482614
rect 516954 482294 517574 482378
rect 516954 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 517574 482294
rect 516954 446614 517574 482058
rect 516954 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 517574 446614
rect 516954 446294 517574 446378
rect 516954 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 517574 446294
rect 516954 410614 517574 446058
rect 516954 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 517574 410614
rect 516954 410294 517574 410378
rect 516954 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 517574 410294
rect 516954 374614 517574 410058
rect 516954 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 517574 374614
rect 516954 374294 517574 374378
rect 516954 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 517574 374294
rect 516954 338614 517574 374058
rect 516954 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 517574 338614
rect 516954 338294 517574 338378
rect 516954 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 517574 338294
rect 516954 302614 517574 338058
rect 516954 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 517574 302614
rect 516954 302294 517574 302378
rect 516954 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 517574 302294
rect 516954 266614 517574 302058
rect 516954 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 517574 266614
rect 516954 266294 517574 266378
rect 516954 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 517574 266294
rect 516954 230614 517574 266058
rect 516954 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 517574 230614
rect 516954 230294 517574 230378
rect 516954 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 517574 230294
rect 516954 194614 517574 230058
rect 516954 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 517574 194614
rect 516954 194294 517574 194378
rect 516954 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 517574 194294
rect 516954 158614 517574 194058
rect 516954 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 517574 158614
rect 516954 158294 517574 158378
rect 516954 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 517574 158294
rect 516954 122614 517574 158058
rect 516954 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 517574 122614
rect 516954 122294 517574 122378
rect 516954 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 517574 122294
rect 516954 86614 517574 122058
rect 516954 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 517574 86614
rect 516954 86294 517574 86378
rect 516954 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 517574 86294
rect 516954 50614 517574 86058
rect 516954 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 517574 50614
rect 516954 50294 517574 50378
rect 516954 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 517574 50294
rect 516954 14614 517574 50058
rect 516954 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 517574 14614
rect 516954 14294 517574 14378
rect 516954 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 517574 14294
rect 498954 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 499574 -7066
rect 498954 -7386 499574 -7302
rect 498954 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 499574 -7386
rect 498954 -7654 499574 -7622
rect 516954 -6106 517574 14058
rect 523794 705798 524414 705830
rect 523794 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 524414 705798
rect 523794 705478 524414 705562
rect 523794 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 524414 705478
rect 523794 669454 524414 705242
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -1306 524414 20898
rect 523794 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 524414 -1306
rect 523794 -1626 524414 -1542
rect 523794 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 524414 -1626
rect 523794 -1894 524414 -1862
rect 527514 673174 528134 707162
rect 527514 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 528134 673174
rect 527514 672854 528134 672938
rect 527514 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 528134 672854
rect 527514 637174 528134 672618
rect 527514 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 528134 637174
rect 527514 636854 528134 636938
rect 527514 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 528134 636854
rect 527514 601174 528134 636618
rect 527514 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 528134 601174
rect 527514 600854 528134 600938
rect 527514 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 528134 600854
rect 527514 565174 528134 600618
rect 527514 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 528134 565174
rect 527514 564854 528134 564938
rect 527514 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 528134 564854
rect 527514 529174 528134 564618
rect 527514 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 528134 529174
rect 527514 528854 528134 528938
rect 527514 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 528134 528854
rect 527514 493174 528134 528618
rect 527514 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 528134 493174
rect 527514 492854 528134 492938
rect 527514 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 528134 492854
rect 527514 457174 528134 492618
rect 527514 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 528134 457174
rect 527514 456854 528134 456938
rect 527514 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 528134 456854
rect 527514 421174 528134 456618
rect 527514 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 528134 421174
rect 527514 420854 528134 420938
rect 527514 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 528134 420854
rect 527514 385174 528134 420618
rect 527514 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 528134 385174
rect 527514 384854 528134 384938
rect 527514 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 528134 384854
rect 527514 349174 528134 384618
rect 527514 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 528134 349174
rect 527514 348854 528134 348938
rect 527514 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 528134 348854
rect 527514 313174 528134 348618
rect 527514 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 528134 313174
rect 527514 312854 528134 312938
rect 527514 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 528134 312854
rect 527514 277174 528134 312618
rect 527514 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 528134 277174
rect 527514 276854 528134 276938
rect 527514 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 528134 276854
rect 527514 241174 528134 276618
rect 527514 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 528134 241174
rect 527514 240854 528134 240938
rect 527514 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 528134 240854
rect 527514 205174 528134 240618
rect 527514 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 528134 205174
rect 527514 204854 528134 204938
rect 527514 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 528134 204854
rect 527514 169174 528134 204618
rect 527514 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 528134 169174
rect 527514 168854 528134 168938
rect 527514 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 528134 168854
rect 527514 133174 528134 168618
rect 527514 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 528134 133174
rect 527514 132854 528134 132938
rect 527514 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 528134 132854
rect 527514 97174 528134 132618
rect 527514 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 528134 97174
rect 527514 96854 528134 96938
rect 527514 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 528134 96854
rect 527514 61174 528134 96618
rect 527514 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 528134 61174
rect 527514 60854 528134 60938
rect 527514 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 528134 60854
rect 527514 25174 528134 60618
rect 527514 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 528134 25174
rect 527514 24854 528134 24938
rect 527514 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 528134 24854
rect 527514 -3226 528134 24618
rect 527514 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 528134 -3226
rect 527514 -3546 528134 -3462
rect 527514 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 528134 -3546
rect 527514 -3814 528134 -3782
rect 531234 676894 531854 709082
rect 531234 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 531854 676894
rect 531234 676574 531854 676658
rect 531234 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 531854 676574
rect 531234 640894 531854 676338
rect 531234 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 531854 640894
rect 531234 640574 531854 640658
rect 531234 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 531854 640574
rect 531234 604894 531854 640338
rect 531234 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 531854 604894
rect 531234 604574 531854 604658
rect 531234 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 531854 604574
rect 531234 568894 531854 604338
rect 531234 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 531854 568894
rect 531234 568574 531854 568658
rect 531234 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 531854 568574
rect 531234 532894 531854 568338
rect 531234 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 531854 532894
rect 531234 532574 531854 532658
rect 531234 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 531854 532574
rect 531234 496894 531854 532338
rect 531234 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 531854 496894
rect 531234 496574 531854 496658
rect 531234 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 531854 496574
rect 531234 460894 531854 496338
rect 531234 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 531854 460894
rect 531234 460574 531854 460658
rect 531234 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 531854 460574
rect 531234 424894 531854 460338
rect 531234 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 531854 424894
rect 531234 424574 531854 424658
rect 531234 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 531854 424574
rect 531234 388894 531854 424338
rect 531234 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 531854 388894
rect 531234 388574 531854 388658
rect 531234 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 531854 388574
rect 531234 352894 531854 388338
rect 531234 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 531854 352894
rect 531234 352574 531854 352658
rect 531234 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 531854 352574
rect 531234 316894 531854 352338
rect 531234 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 531854 316894
rect 531234 316574 531854 316658
rect 531234 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 531854 316574
rect 531234 280894 531854 316338
rect 531234 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 531854 280894
rect 531234 280574 531854 280658
rect 531234 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 531854 280574
rect 531234 244894 531854 280338
rect 531234 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 531854 244894
rect 531234 244574 531854 244658
rect 531234 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 531854 244574
rect 531234 208894 531854 244338
rect 531234 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 531854 208894
rect 531234 208574 531854 208658
rect 531234 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 531854 208574
rect 531234 172894 531854 208338
rect 531234 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 531854 172894
rect 531234 172574 531854 172658
rect 531234 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 531854 172574
rect 531234 136894 531854 172338
rect 531234 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 531854 136894
rect 531234 136574 531854 136658
rect 531234 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 531854 136574
rect 531234 100894 531854 136338
rect 531234 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 531854 100894
rect 531234 100574 531854 100658
rect 531234 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 531854 100574
rect 531234 64894 531854 100338
rect 531234 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 531854 64894
rect 531234 64574 531854 64658
rect 531234 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 531854 64574
rect 531234 28894 531854 64338
rect 531234 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 531854 28894
rect 531234 28574 531854 28658
rect 531234 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 531854 28574
rect 531234 -5146 531854 28338
rect 531234 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 531854 -5146
rect 531234 -5466 531854 -5382
rect 531234 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 531854 -5466
rect 531234 -5734 531854 -5702
rect 534954 680614 535574 711002
rect 552954 710598 553574 711590
rect 552954 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 553574 710598
rect 552954 710278 553574 710362
rect 552954 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 553574 710278
rect 549234 708678 549854 709670
rect 549234 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 549854 708678
rect 549234 708358 549854 708442
rect 549234 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 549854 708358
rect 545514 706758 546134 707750
rect 545514 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 546134 706758
rect 545514 706438 546134 706522
rect 545514 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 546134 706438
rect 534954 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 535574 680614
rect 534954 680294 535574 680378
rect 534954 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 535574 680294
rect 534954 644614 535574 680058
rect 534954 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 535574 644614
rect 534954 644294 535574 644378
rect 534954 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 535574 644294
rect 534954 608614 535574 644058
rect 534954 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 535574 608614
rect 534954 608294 535574 608378
rect 534954 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 535574 608294
rect 534954 572614 535574 608058
rect 534954 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 535574 572614
rect 534954 572294 535574 572378
rect 534954 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 535574 572294
rect 534954 536614 535574 572058
rect 534954 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 535574 536614
rect 534954 536294 535574 536378
rect 534954 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 535574 536294
rect 534954 500614 535574 536058
rect 534954 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 535574 500614
rect 534954 500294 535574 500378
rect 534954 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 535574 500294
rect 534954 464614 535574 500058
rect 534954 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 535574 464614
rect 534954 464294 535574 464378
rect 534954 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 535574 464294
rect 534954 428614 535574 464058
rect 534954 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 535574 428614
rect 534954 428294 535574 428378
rect 534954 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 535574 428294
rect 534954 392614 535574 428058
rect 534954 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 535574 392614
rect 534954 392294 535574 392378
rect 534954 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 535574 392294
rect 534954 356614 535574 392058
rect 534954 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 535574 356614
rect 534954 356294 535574 356378
rect 534954 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 535574 356294
rect 534954 320614 535574 356058
rect 534954 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 535574 320614
rect 534954 320294 535574 320378
rect 534954 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 535574 320294
rect 534954 284614 535574 320058
rect 534954 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 535574 284614
rect 534954 284294 535574 284378
rect 534954 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 535574 284294
rect 534954 248614 535574 284058
rect 534954 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 535574 248614
rect 534954 248294 535574 248378
rect 534954 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 535574 248294
rect 534954 212614 535574 248058
rect 534954 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 535574 212614
rect 534954 212294 535574 212378
rect 534954 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 535574 212294
rect 534954 176614 535574 212058
rect 534954 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 535574 176614
rect 534954 176294 535574 176378
rect 534954 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 535574 176294
rect 534954 140614 535574 176058
rect 534954 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 535574 140614
rect 534954 140294 535574 140378
rect 534954 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 535574 140294
rect 534954 104614 535574 140058
rect 534954 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 535574 104614
rect 534954 104294 535574 104378
rect 534954 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 535574 104294
rect 534954 68614 535574 104058
rect 534954 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 535574 68614
rect 534954 68294 535574 68378
rect 534954 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 535574 68294
rect 534954 32614 535574 68058
rect 534954 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 535574 32614
rect 534954 32294 535574 32378
rect 534954 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 535574 32294
rect 516954 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 517574 -6106
rect 516954 -6426 517574 -6342
rect 516954 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 517574 -6426
rect 516954 -7654 517574 -6662
rect 534954 -7066 535574 32058
rect 541794 704838 542414 705830
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -1894 542414 -902
rect 545514 691174 546134 706202
rect 545514 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 546134 691174
rect 545514 690854 546134 690938
rect 545514 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 546134 690854
rect 545514 655174 546134 690618
rect 545514 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 546134 655174
rect 545514 654854 546134 654938
rect 545514 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 546134 654854
rect 545514 619174 546134 654618
rect 545514 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 546134 619174
rect 545514 618854 546134 618938
rect 545514 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 546134 618854
rect 545514 583174 546134 618618
rect 545514 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 546134 583174
rect 545514 582854 546134 582938
rect 545514 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 546134 582854
rect 545514 547174 546134 582618
rect 545514 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 546134 547174
rect 545514 546854 546134 546938
rect 545514 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 546134 546854
rect 545514 511174 546134 546618
rect 545514 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 546134 511174
rect 545514 510854 546134 510938
rect 545514 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 546134 510854
rect 545514 475174 546134 510618
rect 545514 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 546134 475174
rect 545514 474854 546134 474938
rect 545514 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 546134 474854
rect 545514 439174 546134 474618
rect 545514 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 546134 439174
rect 545514 438854 546134 438938
rect 545514 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 546134 438854
rect 545514 403174 546134 438618
rect 545514 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 546134 403174
rect 545514 402854 546134 402938
rect 545514 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 546134 402854
rect 545514 367174 546134 402618
rect 545514 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 546134 367174
rect 545514 366854 546134 366938
rect 545514 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 546134 366854
rect 545514 331174 546134 366618
rect 545514 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 546134 331174
rect 545514 330854 546134 330938
rect 545514 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 546134 330854
rect 545514 295174 546134 330618
rect 545514 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 546134 295174
rect 545514 294854 546134 294938
rect 545514 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 546134 294854
rect 545514 259174 546134 294618
rect 545514 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 546134 259174
rect 545514 258854 546134 258938
rect 545514 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 546134 258854
rect 545514 223174 546134 258618
rect 545514 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 546134 223174
rect 545514 222854 546134 222938
rect 545514 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 546134 222854
rect 545514 187174 546134 222618
rect 545514 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 546134 187174
rect 545514 186854 546134 186938
rect 545514 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 546134 186854
rect 545514 151174 546134 186618
rect 545514 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 546134 151174
rect 545514 150854 546134 150938
rect 545514 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 546134 150854
rect 545514 115174 546134 150618
rect 545514 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 546134 115174
rect 545514 114854 546134 114938
rect 545514 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 546134 114854
rect 545514 79174 546134 114618
rect 545514 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 546134 79174
rect 545514 78854 546134 78938
rect 545514 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 546134 78854
rect 545514 43174 546134 78618
rect 545514 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 546134 43174
rect 545514 42854 546134 42938
rect 545514 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 546134 42854
rect 545514 7174 546134 42618
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -2266 546134 6618
rect 545514 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 546134 -2266
rect 545514 -2586 546134 -2502
rect 545514 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 546134 -2586
rect 545514 -3814 546134 -2822
rect 549234 694894 549854 708122
rect 549234 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 549854 694894
rect 549234 694574 549854 694658
rect 549234 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 549854 694574
rect 549234 658894 549854 694338
rect 549234 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 549854 658894
rect 549234 658574 549854 658658
rect 549234 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 549854 658574
rect 549234 622894 549854 658338
rect 549234 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 549854 622894
rect 549234 622574 549854 622658
rect 549234 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 549854 622574
rect 549234 586894 549854 622338
rect 549234 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 549854 586894
rect 549234 586574 549854 586658
rect 549234 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 549854 586574
rect 549234 550894 549854 586338
rect 549234 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 549854 550894
rect 549234 550574 549854 550658
rect 549234 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 549854 550574
rect 549234 514894 549854 550338
rect 549234 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 549854 514894
rect 549234 514574 549854 514658
rect 549234 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 549854 514574
rect 549234 478894 549854 514338
rect 549234 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 549854 478894
rect 549234 478574 549854 478658
rect 549234 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 549854 478574
rect 549234 442894 549854 478338
rect 549234 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 549854 442894
rect 549234 442574 549854 442658
rect 549234 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 549854 442574
rect 549234 406894 549854 442338
rect 549234 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 549854 406894
rect 549234 406574 549854 406658
rect 549234 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 549854 406574
rect 549234 370894 549854 406338
rect 549234 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 549854 370894
rect 549234 370574 549854 370658
rect 549234 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 549854 370574
rect 549234 334894 549854 370338
rect 549234 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 549854 334894
rect 549234 334574 549854 334658
rect 549234 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 549854 334574
rect 549234 298894 549854 334338
rect 549234 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 549854 298894
rect 549234 298574 549854 298658
rect 549234 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 549854 298574
rect 549234 262894 549854 298338
rect 549234 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 549854 262894
rect 549234 262574 549854 262658
rect 549234 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 549854 262574
rect 549234 226894 549854 262338
rect 549234 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 549854 226894
rect 549234 226574 549854 226658
rect 549234 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 549854 226574
rect 549234 190894 549854 226338
rect 549234 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 549854 190894
rect 549234 190574 549854 190658
rect 549234 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 549854 190574
rect 549234 154894 549854 190338
rect 549234 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 549854 154894
rect 549234 154574 549854 154658
rect 549234 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 549854 154574
rect 549234 118894 549854 154338
rect 549234 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 549854 118894
rect 549234 118574 549854 118658
rect 549234 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 549854 118574
rect 549234 82894 549854 118338
rect 549234 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 549854 82894
rect 549234 82574 549854 82658
rect 549234 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 549854 82574
rect 549234 46894 549854 82338
rect 549234 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 549854 46894
rect 549234 46574 549854 46658
rect 549234 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 549854 46574
rect 549234 10894 549854 46338
rect 549234 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 549854 10894
rect 549234 10574 549854 10658
rect 549234 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 549854 10574
rect 549234 -4186 549854 10338
rect 549234 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 549854 -4186
rect 549234 -4506 549854 -4422
rect 549234 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 549854 -4506
rect 549234 -5734 549854 -4742
rect 552954 698614 553574 710042
rect 570954 711558 571574 711590
rect 570954 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 571574 711558
rect 570954 711238 571574 711322
rect 570954 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 571574 711238
rect 567234 709638 567854 709670
rect 567234 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 567854 709638
rect 567234 709318 567854 709402
rect 567234 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 567854 709318
rect 563514 707718 564134 707750
rect 563514 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 564134 707718
rect 563514 707398 564134 707482
rect 563514 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 564134 707398
rect 552954 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 553574 698614
rect 552954 698294 553574 698378
rect 552954 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 553574 698294
rect 552954 662614 553574 698058
rect 552954 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 553574 662614
rect 552954 662294 553574 662378
rect 552954 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 553574 662294
rect 552954 626614 553574 662058
rect 552954 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 553574 626614
rect 552954 626294 553574 626378
rect 552954 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 553574 626294
rect 552954 590614 553574 626058
rect 552954 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 553574 590614
rect 552954 590294 553574 590378
rect 552954 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 553574 590294
rect 552954 554614 553574 590058
rect 552954 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 553574 554614
rect 552954 554294 553574 554378
rect 552954 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 553574 554294
rect 552954 518614 553574 554058
rect 552954 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 553574 518614
rect 552954 518294 553574 518378
rect 552954 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 553574 518294
rect 552954 482614 553574 518058
rect 552954 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 553574 482614
rect 552954 482294 553574 482378
rect 552954 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 553574 482294
rect 552954 446614 553574 482058
rect 552954 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 553574 446614
rect 552954 446294 553574 446378
rect 552954 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 553574 446294
rect 552954 410614 553574 446058
rect 552954 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 553574 410614
rect 552954 410294 553574 410378
rect 552954 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 553574 410294
rect 552954 374614 553574 410058
rect 552954 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 553574 374614
rect 552954 374294 553574 374378
rect 552954 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 553574 374294
rect 552954 338614 553574 374058
rect 552954 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 553574 338614
rect 552954 338294 553574 338378
rect 552954 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 553574 338294
rect 552954 302614 553574 338058
rect 552954 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 553574 302614
rect 552954 302294 553574 302378
rect 552954 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 553574 302294
rect 552954 266614 553574 302058
rect 552954 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 553574 266614
rect 552954 266294 553574 266378
rect 552954 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 553574 266294
rect 552954 230614 553574 266058
rect 552954 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 553574 230614
rect 552954 230294 553574 230378
rect 552954 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 553574 230294
rect 552954 194614 553574 230058
rect 552954 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 553574 194614
rect 552954 194294 553574 194378
rect 552954 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 553574 194294
rect 552954 158614 553574 194058
rect 552954 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 553574 158614
rect 552954 158294 553574 158378
rect 552954 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 553574 158294
rect 552954 122614 553574 158058
rect 552954 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 553574 122614
rect 552954 122294 553574 122378
rect 552954 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 553574 122294
rect 552954 86614 553574 122058
rect 552954 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 553574 86614
rect 552954 86294 553574 86378
rect 552954 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 553574 86294
rect 552954 50614 553574 86058
rect 552954 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 553574 50614
rect 552954 50294 553574 50378
rect 552954 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 553574 50294
rect 552954 14614 553574 50058
rect 552954 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 553574 14614
rect 552954 14294 553574 14378
rect 552954 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 553574 14294
rect 534954 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 535574 -7066
rect 534954 -7386 535574 -7302
rect 534954 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 535574 -7386
rect 534954 -7654 535574 -7622
rect 552954 -6106 553574 14058
rect 559794 705798 560414 705830
rect 559794 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 560414 705798
rect 559794 705478 560414 705562
rect 559794 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 560414 705478
rect 559794 669454 560414 705242
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -1306 560414 20898
rect 559794 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 560414 -1306
rect 559794 -1626 560414 -1542
rect 559794 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 560414 -1626
rect 559794 -1894 560414 -1862
rect 563514 673174 564134 707162
rect 563514 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 564134 673174
rect 563514 672854 564134 672938
rect 563514 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 564134 672854
rect 563514 637174 564134 672618
rect 563514 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 564134 637174
rect 563514 636854 564134 636938
rect 563514 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 564134 636854
rect 563514 601174 564134 636618
rect 563514 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 564134 601174
rect 563514 600854 564134 600938
rect 563514 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 564134 600854
rect 563514 565174 564134 600618
rect 563514 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 564134 565174
rect 563514 564854 564134 564938
rect 563514 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 564134 564854
rect 563514 529174 564134 564618
rect 563514 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 564134 529174
rect 563514 528854 564134 528938
rect 563514 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 564134 528854
rect 563514 493174 564134 528618
rect 563514 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 564134 493174
rect 563514 492854 564134 492938
rect 563514 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 564134 492854
rect 563514 457174 564134 492618
rect 563514 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 564134 457174
rect 563514 456854 564134 456938
rect 563514 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 564134 456854
rect 563514 421174 564134 456618
rect 563514 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 564134 421174
rect 563514 420854 564134 420938
rect 563514 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 564134 420854
rect 563514 385174 564134 420618
rect 563514 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 564134 385174
rect 563514 384854 564134 384938
rect 563514 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 564134 384854
rect 563514 349174 564134 384618
rect 563514 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 564134 349174
rect 563514 348854 564134 348938
rect 563514 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 564134 348854
rect 563514 313174 564134 348618
rect 563514 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 564134 313174
rect 563514 312854 564134 312938
rect 563514 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 564134 312854
rect 563514 277174 564134 312618
rect 563514 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 564134 277174
rect 563514 276854 564134 276938
rect 563514 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 564134 276854
rect 563514 241174 564134 276618
rect 563514 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 564134 241174
rect 563514 240854 564134 240938
rect 563514 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 564134 240854
rect 563514 205174 564134 240618
rect 563514 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 564134 205174
rect 563514 204854 564134 204938
rect 563514 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 564134 204854
rect 563514 169174 564134 204618
rect 563514 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 564134 169174
rect 563514 168854 564134 168938
rect 563514 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 564134 168854
rect 563514 133174 564134 168618
rect 563514 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 564134 133174
rect 563514 132854 564134 132938
rect 563514 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 564134 132854
rect 563514 97174 564134 132618
rect 563514 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 564134 97174
rect 563514 96854 564134 96938
rect 563514 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 564134 96854
rect 563514 61174 564134 96618
rect 563514 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 564134 61174
rect 563514 60854 564134 60938
rect 563514 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 564134 60854
rect 563514 25174 564134 60618
rect 563514 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 564134 25174
rect 563514 24854 564134 24938
rect 563514 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 564134 24854
rect 563514 -3226 564134 24618
rect 563514 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 564134 -3226
rect 563514 -3546 564134 -3462
rect 563514 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 564134 -3546
rect 563514 -3814 564134 -3782
rect 567234 676894 567854 709082
rect 567234 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 567854 676894
rect 567234 676574 567854 676658
rect 567234 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 567854 676574
rect 567234 640894 567854 676338
rect 567234 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 567854 640894
rect 567234 640574 567854 640658
rect 567234 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 567854 640574
rect 567234 604894 567854 640338
rect 567234 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 567854 604894
rect 567234 604574 567854 604658
rect 567234 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 567854 604574
rect 567234 568894 567854 604338
rect 567234 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 567854 568894
rect 567234 568574 567854 568658
rect 567234 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 567854 568574
rect 567234 532894 567854 568338
rect 567234 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 567854 532894
rect 567234 532574 567854 532658
rect 567234 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 567854 532574
rect 567234 496894 567854 532338
rect 567234 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 567854 496894
rect 567234 496574 567854 496658
rect 567234 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 567854 496574
rect 567234 460894 567854 496338
rect 567234 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 567854 460894
rect 567234 460574 567854 460658
rect 567234 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 567854 460574
rect 567234 424894 567854 460338
rect 567234 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 567854 424894
rect 567234 424574 567854 424658
rect 567234 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 567854 424574
rect 567234 388894 567854 424338
rect 567234 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 567854 388894
rect 567234 388574 567854 388658
rect 567234 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 567854 388574
rect 567234 352894 567854 388338
rect 567234 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 567854 352894
rect 567234 352574 567854 352658
rect 567234 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 567854 352574
rect 567234 316894 567854 352338
rect 567234 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 567854 316894
rect 567234 316574 567854 316658
rect 567234 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 567854 316574
rect 567234 280894 567854 316338
rect 567234 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 567854 280894
rect 567234 280574 567854 280658
rect 567234 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 567854 280574
rect 567234 244894 567854 280338
rect 567234 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 567854 244894
rect 567234 244574 567854 244658
rect 567234 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 567854 244574
rect 567234 208894 567854 244338
rect 567234 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 567854 208894
rect 567234 208574 567854 208658
rect 567234 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 567854 208574
rect 567234 172894 567854 208338
rect 567234 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 567854 172894
rect 567234 172574 567854 172658
rect 567234 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 567854 172574
rect 567234 136894 567854 172338
rect 567234 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 567854 136894
rect 567234 136574 567854 136658
rect 567234 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 567854 136574
rect 567234 100894 567854 136338
rect 567234 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 567854 100894
rect 567234 100574 567854 100658
rect 567234 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 567854 100574
rect 567234 64894 567854 100338
rect 567234 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 567854 64894
rect 567234 64574 567854 64658
rect 567234 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 567854 64574
rect 567234 28894 567854 64338
rect 567234 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 567854 28894
rect 567234 28574 567854 28658
rect 567234 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 567854 28574
rect 567234 -5146 567854 28338
rect 567234 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 567854 -5146
rect 567234 -5466 567854 -5382
rect 567234 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 567854 -5466
rect 567234 -5734 567854 -5702
rect 570954 680614 571574 711002
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 581514 706758 582134 707750
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 581514 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 582134 706758
rect 581514 706438 582134 706522
rect 581514 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 582134 706438
rect 570954 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 571574 680614
rect 570954 680294 571574 680378
rect 570954 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 571574 680294
rect 570954 644614 571574 680058
rect 570954 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 571574 644614
rect 570954 644294 571574 644378
rect 570954 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 571574 644294
rect 570954 608614 571574 644058
rect 570954 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 571574 608614
rect 570954 608294 571574 608378
rect 570954 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 571574 608294
rect 570954 572614 571574 608058
rect 570954 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 571574 572614
rect 570954 572294 571574 572378
rect 570954 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 571574 572294
rect 570954 536614 571574 572058
rect 570954 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 571574 536614
rect 570954 536294 571574 536378
rect 570954 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 571574 536294
rect 570954 500614 571574 536058
rect 570954 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 571574 500614
rect 570954 500294 571574 500378
rect 570954 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 571574 500294
rect 570954 464614 571574 500058
rect 570954 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 571574 464614
rect 570954 464294 571574 464378
rect 570954 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 571574 464294
rect 570954 428614 571574 464058
rect 570954 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 571574 428614
rect 570954 428294 571574 428378
rect 570954 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 571574 428294
rect 570954 392614 571574 428058
rect 570954 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 571574 392614
rect 570954 392294 571574 392378
rect 570954 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 571574 392294
rect 570954 356614 571574 392058
rect 570954 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 571574 356614
rect 570954 356294 571574 356378
rect 570954 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 571574 356294
rect 570954 320614 571574 356058
rect 570954 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 571574 320614
rect 570954 320294 571574 320378
rect 570954 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 571574 320294
rect 570954 284614 571574 320058
rect 570954 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 571574 284614
rect 570954 284294 571574 284378
rect 570954 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 571574 284294
rect 570954 248614 571574 284058
rect 570954 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 571574 248614
rect 570954 248294 571574 248378
rect 570954 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 571574 248294
rect 570954 212614 571574 248058
rect 570954 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 571574 212614
rect 570954 212294 571574 212378
rect 570954 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 571574 212294
rect 570954 176614 571574 212058
rect 570954 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 571574 176614
rect 570954 176294 571574 176378
rect 570954 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 571574 176294
rect 570954 140614 571574 176058
rect 570954 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 571574 140614
rect 570954 140294 571574 140378
rect 570954 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 571574 140294
rect 570954 104614 571574 140058
rect 570954 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 571574 104614
rect 570954 104294 571574 104378
rect 570954 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 571574 104294
rect 570954 68614 571574 104058
rect 570954 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 571574 68614
rect 570954 68294 571574 68378
rect 570954 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 571574 68294
rect 570954 32614 571574 68058
rect 570954 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 571574 32614
rect 570954 32294 571574 32378
rect 570954 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 571574 32294
rect 552954 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 553574 -6106
rect 552954 -6426 553574 -6342
rect 552954 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 553574 -6426
rect 552954 -7654 553574 -6662
rect 570954 -7066 571574 32058
rect 577794 704838 578414 705830
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 580211 697236 580277 697237
rect 580211 697172 580212 697236
rect 580276 697172 580277 697236
rect 580211 697171 580277 697172
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 580214 177853 580274 697171
rect 581514 691174 582134 706202
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 580395 683908 580461 683909
rect 580395 683844 580396 683908
rect 580460 683844 580461 683908
rect 580395 683843 580461 683844
rect 580398 179621 580458 683843
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 580395 179620 580461 179621
rect 580395 179556 580396 179620
rect 580460 179556 580461 179620
rect 580395 179555 580461 179556
rect 580211 177852 580277 177853
rect 580211 177788 580212 177852
rect 580276 177788 580277 177852
rect 580211 177787 580277 177788
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -1894 578414 -902
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -2266 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 669454 586890 705242
rect 586270 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect 586270 669134 586890 669218
rect 586270 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect 586270 633454 586890 668898
rect 586270 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect 586270 633134 586890 633218
rect 586270 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect 586270 597454 586890 632898
rect 586270 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect 586270 597134 586890 597218
rect 586270 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect 586270 561454 586890 596898
rect 586270 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect 586270 561134 586890 561218
rect 586270 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect 586270 525454 586890 560898
rect 586270 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect 586270 525134 586890 525218
rect 586270 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect 586270 489454 586890 524898
rect 586270 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect 586270 489134 586890 489218
rect 586270 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect 586270 453454 586890 488898
rect 586270 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect 586270 453134 586890 453218
rect 586270 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect 586270 417454 586890 452898
rect 586270 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect 586270 417134 586890 417218
rect 586270 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect 586270 381454 586890 416898
rect 586270 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect 586270 381134 586890 381218
rect 586270 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect 586270 345454 586890 380898
rect 586270 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect 586270 345134 586890 345218
rect 586270 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect 586270 309454 586890 344898
rect 586270 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect 586270 309134 586890 309218
rect 586270 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect 586270 273454 586890 308898
rect 586270 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect 586270 273134 586890 273218
rect 586270 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect 586270 237454 586890 272898
rect 586270 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect 586270 237134 586890 237218
rect 586270 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect 586270 201454 586890 236898
rect 586270 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect 586270 201134 586890 201218
rect 586270 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect 586270 165454 586890 200898
rect 586270 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect 586270 165134 586890 165218
rect 586270 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect 586270 129454 586890 164898
rect 586270 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect 586270 129134 586890 129218
rect 586270 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect 586270 93454 586890 128898
rect 586270 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect 586270 93134 586890 93218
rect 586270 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect 586270 57454 586890 92898
rect 586270 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect 586270 57134 586890 57218
rect 586270 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect 586270 21454 586890 56898
rect 586270 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect 586270 21134 586890 21218
rect 586270 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect 586270 -1306 586890 20898
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 691174 587850 706202
rect 587230 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 587850 691174
rect 587230 690854 587850 690938
rect 587230 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 587850 690854
rect 587230 655174 587850 690618
rect 587230 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 587850 655174
rect 587230 654854 587850 654938
rect 587230 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 587850 654854
rect 587230 619174 587850 654618
rect 587230 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 587850 619174
rect 587230 618854 587850 618938
rect 587230 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 587850 618854
rect 587230 583174 587850 618618
rect 587230 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 587850 583174
rect 587230 582854 587850 582938
rect 587230 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 587850 582854
rect 587230 547174 587850 582618
rect 587230 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 587850 547174
rect 587230 546854 587850 546938
rect 587230 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 587850 546854
rect 587230 511174 587850 546618
rect 587230 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 587850 511174
rect 587230 510854 587850 510938
rect 587230 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 587850 510854
rect 587230 475174 587850 510618
rect 587230 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 587850 475174
rect 587230 474854 587850 474938
rect 587230 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 587850 474854
rect 587230 439174 587850 474618
rect 587230 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 587850 439174
rect 587230 438854 587850 438938
rect 587230 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 587850 438854
rect 587230 403174 587850 438618
rect 587230 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 587850 403174
rect 587230 402854 587850 402938
rect 587230 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 587850 402854
rect 587230 367174 587850 402618
rect 587230 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 587850 367174
rect 587230 366854 587850 366938
rect 587230 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 587850 366854
rect 587230 331174 587850 366618
rect 587230 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 587850 331174
rect 587230 330854 587850 330938
rect 587230 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 587850 330854
rect 587230 295174 587850 330618
rect 587230 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 587850 295174
rect 587230 294854 587850 294938
rect 587230 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 587850 294854
rect 587230 259174 587850 294618
rect 587230 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 587850 259174
rect 587230 258854 587850 258938
rect 587230 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 587850 258854
rect 587230 223174 587850 258618
rect 587230 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 587850 223174
rect 587230 222854 587850 222938
rect 587230 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 587850 222854
rect 587230 187174 587850 222618
rect 587230 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 587850 187174
rect 587230 186854 587850 186938
rect 587230 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 587850 186854
rect 587230 151174 587850 186618
rect 587230 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 587850 151174
rect 587230 150854 587850 150938
rect 587230 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 587850 150854
rect 587230 115174 587850 150618
rect 587230 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 587850 115174
rect 587230 114854 587850 114938
rect 587230 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 587850 114854
rect 587230 79174 587850 114618
rect 587230 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 587850 79174
rect 587230 78854 587850 78938
rect 587230 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 587850 78854
rect 587230 43174 587850 78618
rect 587230 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 587850 43174
rect 587230 42854 587850 42938
rect 587230 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 587850 42854
rect 587230 7174 587850 42618
rect 587230 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 587850 7174
rect 587230 6854 587850 6938
rect 587230 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 587850 6854
rect 581514 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 582134 -2266
rect 581514 -2586 582134 -2502
rect 581514 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 582134 -2586
rect 581514 -3814 582134 -2822
rect 587230 -2266 587850 6618
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 673174 588810 707162
rect 588190 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect 588190 672854 588810 672938
rect 588190 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect 588190 637174 588810 672618
rect 588190 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect 588190 636854 588810 636938
rect 588190 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect 588190 601174 588810 636618
rect 588190 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect 588190 600854 588810 600938
rect 588190 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect 588190 565174 588810 600618
rect 588190 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect 588190 564854 588810 564938
rect 588190 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect 588190 529174 588810 564618
rect 588190 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect 588190 528854 588810 528938
rect 588190 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect 588190 493174 588810 528618
rect 588190 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect 588190 492854 588810 492938
rect 588190 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect 588190 457174 588810 492618
rect 588190 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect 588190 456854 588810 456938
rect 588190 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect 588190 421174 588810 456618
rect 588190 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect 588190 420854 588810 420938
rect 588190 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect 588190 385174 588810 420618
rect 588190 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect 588190 384854 588810 384938
rect 588190 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect 588190 349174 588810 384618
rect 588190 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect 588190 348854 588810 348938
rect 588190 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect 588190 313174 588810 348618
rect 588190 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect 588190 312854 588810 312938
rect 588190 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect 588190 277174 588810 312618
rect 588190 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect 588190 276854 588810 276938
rect 588190 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect 588190 241174 588810 276618
rect 588190 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect 588190 240854 588810 240938
rect 588190 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect 588190 205174 588810 240618
rect 588190 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect 588190 204854 588810 204938
rect 588190 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect 588190 169174 588810 204618
rect 588190 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect 588190 168854 588810 168938
rect 588190 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect 588190 133174 588810 168618
rect 588190 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect 588190 132854 588810 132938
rect 588190 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect 588190 97174 588810 132618
rect 588190 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect 588190 96854 588810 96938
rect 588190 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect 588190 61174 588810 96618
rect 588190 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect 588190 60854 588810 60938
rect 588190 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect 588190 25174 588810 60618
rect 588190 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect 588190 24854 588810 24938
rect 588190 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect 588190 -3226 588810 24618
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 694894 589770 708122
rect 589150 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 589770 694894
rect 589150 694574 589770 694658
rect 589150 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 589770 694574
rect 589150 658894 589770 694338
rect 589150 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 589770 658894
rect 589150 658574 589770 658658
rect 589150 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 589770 658574
rect 589150 622894 589770 658338
rect 589150 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 589770 622894
rect 589150 622574 589770 622658
rect 589150 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 589770 622574
rect 589150 586894 589770 622338
rect 589150 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 589770 586894
rect 589150 586574 589770 586658
rect 589150 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 589770 586574
rect 589150 550894 589770 586338
rect 589150 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 589770 550894
rect 589150 550574 589770 550658
rect 589150 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 589770 550574
rect 589150 514894 589770 550338
rect 589150 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 589770 514894
rect 589150 514574 589770 514658
rect 589150 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 589770 514574
rect 589150 478894 589770 514338
rect 589150 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 589770 478894
rect 589150 478574 589770 478658
rect 589150 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 589770 478574
rect 589150 442894 589770 478338
rect 589150 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 589770 442894
rect 589150 442574 589770 442658
rect 589150 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 589770 442574
rect 589150 406894 589770 442338
rect 589150 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 589770 406894
rect 589150 406574 589770 406658
rect 589150 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 589770 406574
rect 589150 370894 589770 406338
rect 589150 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 589770 370894
rect 589150 370574 589770 370658
rect 589150 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 589770 370574
rect 589150 334894 589770 370338
rect 589150 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 589770 334894
rect 589150 334574 589770 334658
rect 589150 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 589770 334574
rect 589150 298894 589770 334338
rect 589150 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 589770 298894
rect 589150 298574 589770 298658
rect 589150 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 589770 298574
rect 589150 262894 589770 298338
rect 589150 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 589770 262894
rect 589150 262574 589770 262658
rect 589150 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 589770 262574
rect 589150 226894 589770 262338
rect 589150 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 589770 226894
rect 589150 226574 589770 226658
rect 589150 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 589770 226574
rect 589150 190894 589770 226338
rect 589150 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 589770 190894
rect 589150 190574 589770 190658
rect 589150 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 589770 190574
rect 589150 154894 589770 190338
rect 589150 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 589770 154894
rect 589150 154574 589770 154658
rect 589150 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 589770 154574
rect 589150 118894 589770 154338
rect 589150 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 589770 118894
rect 589150 118574 589770 118658
rect 589150 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 589770 118574
rect 589150 82894 589770 118338
rect 589150 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 589770 82894
rect 589150 82574 589770 82658
rect 589150 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 589770 82574
rect 589150 46894 589770 82338
rect 589150 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 589770 46894
rect 589150 46574 589770 46658
rect 589150 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 589770 46574
rect 589150 10894 589770 46338
rect 589150 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 589770 10894
rect 589150 10574 589770 10658
rect 589150 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 589770 10574
rect 589150 -4186 589770 10338
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 676894 590730 709082
rect 590110 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect 590110 676574 590730 676658
rect 590110 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect 590110 640894 590730 676338
rect 590110 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect 590110 640574 590730 640658
rect 590110 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect 590110 604894 590730 640338
rect 590110 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect 590110 604574 590730 604658
rect 590110 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect 590110 568894 590730 604338
rect 590110 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect 590110 568574 590730 568658
rect 590110 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect 590110 532894 590730 568338
rect 590110 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect 590110 532574 590730 532658
rect 590110 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect 590110 496894 590730 532338
rect 590110 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect 590110 496574 590730 496658
rect 590110 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect 590110 460894 590730 496338
rect 590110 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect 590110 460574 590730 460658
rect 590110 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect 590110 424894 590730 460338
rect 590110 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect 590110 424574 590730 424658
rect 590110 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect 590110 388894 590730 424338
rect 590110 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect 590110 388574 590730 388658
rect 590110 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect 590110 352894 590730 388338
rect 590110 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect 590110 352574 590730 352658
rect 590110 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect 590110 316894 590730 352338
rect 590110 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect 590110 316574 590730 316658
rect 590110 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect 590110 280894 590730 316338
rect 590110 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect 590110 280574 590730 280658
rect 590110 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect 590110 244894 590730 280338
rect 590110 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect 590110 244574 590730 244658
rect 590110 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect 590110 208894 590730 244338
rect 590110 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect 590110 208574 590730 208658
rect 590110 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect 590110 172894 590730 208338
rect 590110 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect 590110 172574 590730 172658
rect 590110 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect 590110 136894 590730 172338
rect 590110 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect 590110 136574 590730 136658
rect 590110 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect 590110 100894 590730 136338
rect 590110 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect 590110 100574 590730 100658
rect 590110 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect 590110 64894 590730 100338
rect 590110 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect 590110 64574 590730 64658
rect 590110 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect 590110 28894 590730 64338
rect 590110 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect 590110 28574 590730 28658
rect 590110 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect 590110 -5146 590730 28338
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 698614 591690 710042
rect 591070 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 591690 698614
rect 591070 698294 591690 698378
rect 591070 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 591690 698294
rect 591070 662614 591690 698058
rect 591070 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 591690 662614
rect 591070 662294 591690 662378
rect 591070 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 591690 662294
rect 591070 626614 591690 662058
rect 591070 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 591690 626614
rect 591070 626294 591690 626378
rect 591070 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 591690 626294
rect 591070 590614 591690 626058
rect 591070 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 591690 590614
rect 591070 590294 591690 590378
rect 591070 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 591690 590294
rect 591070 554614 591690 590058
rect 591070 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 591690 554614
rect 591070 554294 591690 554378
rect 591070 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 591690 554294
rect 591070 518614 591690 554058
rect 591070 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 591690 518614
rect 591070 518294 591690 518378
rect 591070 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 591690 518294
rect 591070 482614 591690 518058
rect 591070 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 591690 482614
rect 591070 482294 591690 482378
rect 591070 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 591690 482294
rect 591070 446614 591690 482058
rect 591070 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 591690 446614
rect 591070 446294 591690 446378
rect 591070 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 591690 446294
rect 591070 410614 591690 446058
rect 591070 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 591690 410614
rect 591070 410294 591690 410378
rect 591070 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 591690 410294
rect 591070 374614 591690 410058
rect 591070 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 591690 374614
rect 591070 374294 591690 374378
rect 591070 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 591690 374294
rect 591070 338614 591690 374058
rect 591070 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 591690 338614
rect 591070 338294 591690 338378
rect 591070 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 591690 338294
rect 591070 302614 591690 338058
rect 591070 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 591690 302614
rect 591070 302294 591690 302378
rect 591070 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 591690 302294
rect 591070 266614 591690 302058
rect 591070 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 591690 266614
rect 591070 266294 591690 266378
rect 591070 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 591690 266294
rect 591070 230614 591690 266058
rect 591070 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 591690 230614
rect 591070 230294 591690 230378
rect 591070 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 591690 230294
rect 591070 194614 591690 230058
rect 591070 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 591690 194614
rect 591070 194294 591690 194378
rect 591070 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 591690 194294
rect 591070 158614 591690 194058
rect 591070 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 591690 158614
rect 591070 158294 591690 158378
rect 591070 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 591690 158294
rect 591070 122614 591690 158058
rect 591070 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 591690 122614
rect 591070 122294 591690 122378
rect 591070 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 591690 122294
rect 591070 86614 591690 122058
rect 591070 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 591690 86614
rect 591070 86294 591690 86378
rect 591070 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 591690 86294
rect 591070 50614 591690 86058
rect 591070 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 591690 50614
rect 591070 50294 591690 50378
rect 591070 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 591690 50294
rect 591070 14614 591690 50058
rect 591070 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 591690 14614
rect 591070 14294 591690 14378
rect 591070 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 591690 14294
rect 591070 -6106 591690 14058
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 680614 592650 711002
rect 592030 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect 592030 680294 592650 680378
rect 592030 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect 592030 644614 592650 680058
rect 592030 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect 592030 644294 592650 644378
rect 592030 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect 592030 608614 592650 644058
rect 592030 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect 592030 608294 592650 608378
rect 592030 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect 592030 572614 592650 608058
rect 592030 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect 592030 572294 592650 572378
rect 592030 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect 592030 536614 592650 572058
rect 592030 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect 592030 536294 592650 536378
rect 592030 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect 592030 500614 592650 536058
rect 592030 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect 592030 500294 592650 500378
rect 592030 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect 592030 464614 592650 500058
rect 592030 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect 592030 464294 592650 464378
rect 592030 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect 592030 428614 592650 464058
rect 592030 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect 592030 428294 592650 428378
rect 592030 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect 592030 392614 592650 428058
rect 592030 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect 592030 392294 592650 392378
rect 592030 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect 592030 356614 592650 392058
rect 592030 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect 592030 356294 592650 356378
rect 592030 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect 592030 320614 592650 356058
rect 592030 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect 592030 320294 592650 320378
rect 592030 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect 592030 284614 592650 320058
rect 592030 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect 592030 284294 592650 284378
rect 592030 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect 592030 248614 592650 284058
rect 592030 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect 592030 248294 592650 248378
rect 592030 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect 592030 212614 592650 248058
rect 592030 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect 592030 212294 592650 212378
rect 592030 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect 592030 176614 592650 212058
rect 592030 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect 592030 176294 592650 176378
rect 592030 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect 592030 140614 592650 176058
rect 592030 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect 592030 140294 592650 140378
rect 592030 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect 592030 104614 592650 140058
rect 592030 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect 592030 104294 592650 104378
rect 592030 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect 592030 68614 592650 104058
rect 592030 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect 592030 68294 592650 68378
rect 592030 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect 592030 32614 592650 68058
rect 592030 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect 592030 32294 592650 32378
rect 592030 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect 570954 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 571574 -7066
rect 570954 -7386 571574 -7302
rect 570954 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 571574 -7386
rect 570954 -7654 571574 -7622
rect 592030 -7066 592650 32058
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 680378 -8458 680614
rect -8374 680378 -8138 680614
rect -8694 680058 -8458 680294
rect -8374 680058 -8138 680294
rect -8694 644378 -8458 644614
rect -8374 644378 -8138 644614
rect -8694 644058 -8458 644294
rect -8374 644058 -8138 644294
rect -8694 608378 -8458 608614
rect -8374 608378 -8138 608614
rect -8694 608058 -8458 608294
rect -8374 608058 -8138 608294
rect -8694 572378 -8458 572614
rect -8374 572378 -8138 572614
rect -8694 572058 -8458 572294
rect -8374 572058 -8138 572294
rect -8694 536378 -8458 536614
rect -8374 536378 -8138 536614
rect -8694 536058 -8458 536294
rect -8374 536058 -8138 536294
rect -8694 500378 -8458 500614
rect -8374 500378 -8138 500614
rect -8694 500058 -8458 500294
rect -8374 500058 -8138 500294
rect -8694 464378 -8458 464614
rect -8374 464378 -8138 464614
rect -8694 464058 -8458 464294
rect -8374 464058 -8138 464294
rect -8694 428378 -8458 428614
rect -8374 428378 -8138 428614
rect -8694 428058 -8458 428294
rect -8374 428058 -8138 428294
rect -8694 392378 -8458 392614
rect -8374 392378 -8138 392614
rect -8694 392058 -8458 392294
rect -8374 392058 -8138 392294
rect -8694 356378 -8458 356614
rect -8374 356378 -8138 356614
rect -8694 356058 -8458 356294
rect -8374 356058 -8138 356294
rect -8694 320378 -8458 320614
rect -8374 320378 -8138 320614
rect -8694 320058 -8458 320294
rect -8374 320058 -8138 320294
rect -8694 284378 -8458 284614
rect -8374 284378 -8138 284614
rect -8694 284058 -8458 284294
rect -8374 284058 -8138 284294
rect -8694 248378 -8458 248614
rect -8374 248378 -8138 248614
rect -8694 248058 -8458 248294
rect -8374 248058 -8138 248294
rect -8694 212378 -8458 212614
rect -8374 212378 -8138 212614
rect -8694 212058 -8458 212294
rect -8374 212058 -8138 212294
rect -8694 176378 -8458 176614
rect -8374 176378 -8138 176614
rect -8694 176058 -8458 176294
rect -8374 176058 -8138 176294
rect -8694 140378 -8458 140614
rect -8374 140378 -8138 140614
rect -8694 140058 -8458 140294
rect -8374 140058 -8138 140294
rect -8694 104378 -8458 104614
rect -8374 104378 -8138 104614
rect -8694 104058 -8458 104294
rect -8374 104058 -8138 104294
rect -8694 68378 -8458 68614
rect -8374 68378 -8138 68614
rect -8694 68058 -8458 68294
rect -8374 68058 -8138 68294
rect -8694 32378 -8458 32614
rect -8374 32378 -8138 32614
rect -8694 32058 -8458 32294
rect -8374 32058 -8138 32294
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect 12986 710362 13222 710598
rect 13306 710362 13542 710598
rect 12986 710042 13222 710278
rect 13306 710042 13542 710278
rect -7734 698378 -7498 698614
rect -7414 698378 -7178 698614
rect -7734 698058 -7498 698294
rect -7414 698058 -7178 698294
rect -7734 662378 -7498 662614
rect -7414 662378 -7178 662614
rect -7734 662058 -7498 662294
rect -7414 662058 -7178 662294
rect -7734 626378 -7498 626614
rect -7414 626378 -7178 626614
rect -7734 626058 -7498 626294
rect -7414 626058 -7178 626294
rect -7734 590378 -7498 590614
rect -7414 590378 -7178 590614
rect -7734 590058 -7498 590294
rect -7414 590058 -7178 590294
rect -7734 554378 -7498 554614
rect -7414 554378 -7178 554614
rect -7734 554058 -7498 554294
rect -7414 554058 -7178 554294
rect -7734 518378 -7498 518614
rect -7414 518378 -7178 518614
rect -7734 518058 -7498 518294
rect -7414 518058 -7178 518294
rect -7734 482378 -7498 482614
rect -7414 482378 -7178 482614
rect -7734 482058 -7498 482294
rect -7414 482058 -7178 482294
rect -7734 446378 -7498 446614
rect -7414 446378 -7178 446614
rect -7734 446058 -7498 446294
rect -7414 446058 -7178 446294
rect -7734 410378 -7498 410614
rect -7414 410378 -7178 410614
rect -7734 410058 -7498 410294
rect -7414 410058 -7178 410294
rect -7734 374378 -7498 374614
rect -7414 374378 -7178 374614
rect -7734 374058 -7498 374294
rect -7414 374058 -7178 374294
rect -7734 338378 -7498 338614
rect -7414 338378 -7178 338614
rect -7734 338058 -7498 338294
rect -7414 338058 -7178 338294
rect -7734 302378 -7498 302614
rect -7414 302378 -7178 302614
rect -7734 302058 -7498 302294
rect -7414 302058 -7178 302294
rect -7734 266378 -7498 266614
rect -7414 266378 -7178 266614
rect -7734 266058 -7498 266294
rect -7414 266058 -7178 266294
rect -7734 230378 -7498 230614
rect -7414 230378 -7178 230614
rect -7734 230058 -7498 230294
rect -7414 230058 -7178 230294
rect -7734 194378 -7498 194614
rect -7414 194378 -7178 194614
rect -7734 194058 -7498 194294
rect -7414 194058 -7178 194294
rect -7734 158378 -7498 158614
rect -7414 158378 -7178 158614
rect -7734 158058 -7498 158294
rect -7414 158058 -7178 158294
rect -7734 122378 -7498 122614
rect -7414 122378 -7178 122614
rect -7734 122058 -7498 122294
rect -7414 122058 -7178 122294
rect -7734 86378 -7498 86614
rect -7414 86378 -7178 86614
rect -7734 86058 -7498 86294
rect -7414 86058 -7178 86294
rect -7734 50378 -7498 50614
rect -7414 50378 -7178 50614
rect -7734 50058 -7498 50294
rect -7414 50058 -7178 50294
rect -7734 14378 -7498 14614
rect -7414 14378 -7178 14614
rect -7734 14058 -7498 14294
rect -7414 14058 -7178 14294
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 676658 -6538 676894
rect -6454 676658 -6218 676894
rect -6774 676338 -6538 676574
rect -6454 676338 -6218 676574
rect -6774 640658 -6538 640894
rect -6454 640658 -6218 640894
rect -6774 640338 -6538 640574
rect -6454 640338 -6218 640574
rect -6774 604658 -6538 604894
rect -6454 604658 -6218 604894
rect -6774 604338 -6538 604574
rect -6454 604338 -6218 604574
rect -6774 568658 -6538 568894
rect -6454 568658 -6218 568894
rect -6774 568338 -6538 568574
rect -6454 568338 -6218 568574
rect -6774 532658 -6538 532894
rect -6454 532658 -6218 532894
rect -6774 532338 -6538 532574
rect -6454 532338 -6218 532574
rect -6774 496658 -6538 496894
rect -6454 496658 -6218 496894
rect -6774 496338 -6538 496574
rect -6454 496338 -6218 496574
rect -6774 460658 -6538 460894
rect -6454 460658 -6218 460894
rect -6774 460338 -6538 460574
rect -6454 460338 -6218 460574
rect -6774 424658 -6538 424894
rect -6454 424658 -6218 424894
rect -6774 424338 -6538 424574
rect -6454 424338 -6218 424574
rect -6774 388658 -6538 388894
rect -6454 388658 -6218 388894
rect -6774 388338 -6538 388574
rect -6454 388338 -6218 388574
rect -6774 352658 -6538 352894
rect -6454 352658 -6218 352894
rect -6774 352338 -6538 352574
rect -6454 352338 -6218 352574
rect -6774 316658 -6538 316894
rect -6454 316658 -6218 316894
rect -6774 316338 -6538 316574
rect -6454 316338 -6218 316574
rect -6774 280658 -6538 280894
rect -6454 280658 -6218 280894
rect -6774 280338 -6538 280574
rect -6454 280338 -6218 280574
rect -6774 244658 -6538 244894
rect -6454 244658 -6218 244894
rect -6774 244338 -6538 244574
rect -6454 244338 -6218 244574
rect -6774 208658 -6538 208894
rect -6454 208658 -6218 208894
rect -6774 208338 -6538 208574
rect -6454 208338 -6218 208574
rect -6774 172658 -6538 172894
rect -6454 172658 -6218 172894
rect -6774 172338 -6538 172574
rect -6454 172338 -6218 172574
rect -6774 136658 -6538 136894
rect -6454 136658 -6218 136894
rect -6774 136338 -6538 136574
rect -6454 136338 -6218 136574
rect -6774 100658 -6538 100894
rect -6454 100658 -6218 100894
rect -6774 100338 -6538 100574
rect -6454 100338 -6218 100574
rect -6774 64658 -6538 64894
rect -6454 64658 -6218 64894
rect -6774 64338 -6538 64574
rect -6454 64338 -6218 64574
rect -6774 28658 -6538 28894
rect -6454 28658 -6218 28894
rect -6774 28338 -6538 28574
rect -6454 28338 -6218 28574
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect 9266 708442 9502 708678
rect 9586 708442 9822 708678
rect 9266 708122 9502 708358
rect 9586 708122 9822 708358
rect -5814 694658 -5578 694894
rect -5494 694658 -5258 694894
rect -5814 694338 -5578 694574
rect -5494 694338 -5258 694574
rect -5814 658658 -5578 658894
rect -5494 658658 -5258 658894
rect -5814 658338 -5578 658574
rect -5494 658338 -5258 658574
rect -5814 622658 -5578 622894
rect -5494 622658 -5258 622894
rect -5814 622338 -5578 622574
rect -5494 622338 -5258 622574
rect -5814 586658 -5578 586894
rect -5494 586658 -5258 586894
rect -5814 586338 -5578 586574
rect -5494 586338 -5258 586574
rect -5814 550658 -5578 550894
rect -5494 550658 -5258 550894
rect -5814 550338 -5578 550574
rect -5494 550338 -5258 550574
rect -5814 514658 -5578 514894
rect -5494 514658 -5258 514894
rect -5814 514338 -5578 514574
rect -5494 514338 -5258 514574
rect -5814 478658 -5578 478894
rect -5494 478658 -5258 478894
rect -5814 478338 -5578 478574
rect -5494 478338 -5258 478574
rect -5814 442658 -5578 442894
rect -5494 442658 -5258 442894
rect -5814 442338 -5578 442574
rect -5494 442338 -5258 442574
rect -5814 406658 -5578 406894
rect -5494 406658 -5258 406894
rect -5814 406338 -5578 406574
rect -5494 406338 -5258 406574
rect -5814 370658 -5578 370894
rect -5494 370658 -5258 370894
rect -5814 370338 -5578 370574
rect -5494 370338 -5258 370574
rect -5814 334658 -5578 334894
rect -5494 334658 -5258 334894
rect -5814 334338 -5578 334574
rect -5494 334338 -5258 334574
rect -5814 298658 -5578 298894
rect -5494 298658 -5258 298894
rect -5814 298338 -5578 298574
rect -5494 298338 -5258 298574
rect -5814 262658 -5578 262894
rect -5494 262658 -5258 262894
rect -5814 262338 -5578 262574
rect -5494 262338 -5258 262574
rect -5814 226658 -5578 226894
rect -5494 226658 -5258 226894
rect -5814 226338 -5578 226574
rect -5494 226338 -5258 226574
rect -5814 190658 -5578 190894
rect -5494 190658 -5258 190894
rect -5814 190338 -5578 190574
rect -5494 190338 -5258 190574
rect -5814 154658 -5578 154894
rect -5494 154658 -5258 154894
rect -5814 154338 -5578 154574
rect -5494 154338 -5258 154574
rect -5814 118658 -5578 118894
rect -5494 118658 -5258 118894
rect -5814 118338 -5578 118574
rect -5494 118338 -5258 118574
rect -5814 82658 -5578 82894
rect -5494 82658 -5258 82894
rect -5814 82338 -5578 82574
rect -5494 82338 -5258 82574
rect -5814 46658 -5578 46894
rect -5494 46658 -5258 46894
rect -5814 46338 -5578 46574
rect -5494 46338 -5258 46574
rect -5814 10658 -5578 10894
rect -5494 10658 -5258 10894
rect -5814 10338 -5578 10574
rect -5494 10338 -5258 10574
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 672938 -4618 673174
rect -4534 672938 -4298 673174
rect -4854 672618 -4618 672854
rect -4534 672618 -4298 672854
rect -4854 636938 -4618 637174
rect -4534 636938 -4298 637174
rect -4854 636618 -4618 636854
rect -4534 636618 -4298 636854
rect -4854 600938 -4618 601174
rect -4534 600938 -4298 601174
rect -4854 600618 -4618 600854
rect -4534 600618 -4298 600854
rect -4854 564938 -4618 565174
rect -4534 564938 -4298 565174
rect -4854 564618 -4618 564854
rect -4534 564618 -4298 564854
rect -4854 528938 -4618 529174
rect -4534 528938 -4298 529174
rect -4854 528618 -4618 528854
rect -4534 528618 -4298 528854
rect -4854 492938 -4618 493174
rect -4534 492938 -4298 493174
rect -4854 492618 -4618 492854
rect -4534 492618 -4298 492854
rect -4854 456938 -4618 457174
rect -4534 456938 -4298 457174
rect -4854 456618 -4618 456854
rect -4534 456618 -4298 456854
rect -4854 420938 -4618 421174
rect -4534 420938 -4298 421174
rect -4854 420618 -4618 420854
rect -4534 420618 -4298 420854
rect -4854 384938 -4618 385174
rect -4534 384938 -4298 385174
rect -4854 384618 -4618 384854
rect -4534 384618 -4298 384854
rect -4854 348938 -4618 349174
rect -4534 348938 -4298 349174
rect -4854 348618 -4618 348854
rect -4534 348618 -4298 348854
rect -4854 312938 -4618 313174
rect -4534 312938 -4298 313174
rect -4854 312618 -4618 312854
rect -4534 312618 -4298 312854
rect -4854 276938 -4618 277174
rect -4534 276938 -4298 277174
rect -4854 276618 -4618 276854
rect -4534 276618 -4298 276854
rect -4854 240938 -4618 241174
rect -4534 240938 -4298 241174
rect -4854 240618 -4618 240854
rect -4534 240618 -4298 240854
rect -4854 204938 -4618 205174
rect -4534 204938 -4298 205174
rect -4854 204618 -4618 204854
rect -4534 204618 -4298 204854
rect -4854 168938 -4618 169174
rect -4534 168938 -4298 169174
rect -4854 168618 -4618 168854
rect -4534 168618 -4298 168854
rect -4854 132938 -4618 133174
rect -4534 132938 -4298 133174
rect -4854 132618 -4618 132854
rect -4534 132618 -4298 132854
rect -4854 96938 -4618 97174
rect -4534 96938 -4298 97174
rect -4854 96618 -4618 96854
rect -4534 96618 -4298 96854
rect -4854 60938 -4618 61174
rect -4534 60938 -4298 61174
rect -4854 60618 -4618 60854
rect -4534 60618 -4298 60854
rect -4854 24938 -4618 25174
rect -4534 24938 -4298 25174
rect -4854 24618 -4618 24854
rect -4534 24618 -4298 24854
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect 5546 706522 5782 706758
rect 5866 706522 6102 706758
rect 5546 706202 5782 706438
rect 5866 706202 6102 706438
rect -3894 690938 -3658 691174
rect -3574 690938 -3338 691174
rect -3894 690618 -3658 690854
rect -3574 690618 -3338 690854
rect -3894 654938 -3658 655174
rect -3574 654938 -3338 655174
rect -3894 654618 -3658 654854
rect -3574 654618 -3338 654854
rect -3894 618938 -3658 619174
rect -3574 618938 -3338 619174
rect -3894 618618 -3658 618854
rect -3574 618618 -3338 618854
rect -3894 582938 -3658 583174
rect -3574 582938 -3338 583174
rect -3894 582618 -3658 582854
rect -3574 582618 -3338 582854
rect -3894 546938 -3658 547174
rect -3574 546938 -3338 547174
rect -3894 546618 -3658 546854
rect -3574 546618 -3338 546854
rect -3894 510938 -3658 511174
rect -3574 510938 -3338 511174
rect -3894 510618 -3658 510854
rect -3574 510618 -3338 510854
rect -3894 474938 -3658 475174
rect -3574 474938 -3338 475174
rect -3894 474618 -3658 474854
rect -3574 474618 -3338 474854
rect -3894 438938 -3658 439174
rect -3574 438938 -3338 439174
rect -3894 438618 -3658 438854
rect -3574 438618 -3338 438854
rect -3894 402938 -3658 403174
rect -3574 402938 -3338 403174
rect -3894 402618 -3658 402854
rect -3574 402618 -3338 402854
rect -3894 366938 -3658 367174
rect -3574 366938 -3338 367174
rect -3894 366618 -3658 366854
rect -3574 366618 -3338 366854
rect -3894 330938 -3658 331174
rect -3574 330938 -3338 331174
rect -3894 330618 -3658 330854
rect -3574 330618 -3338 330854
rect -3894 294938 -3658 295174
rect -3574 294938 -3338 295174
rect -3894 294618 -3658 294854
rect -3574 294618 -3338 294854
rect -3894 258938 -3658 259174
rect -3574 258938 -3338 259174
rect -3894 258618 -3658 258854
rect -3574 258618 -3338 258854
rect -3894 222938 -3658 223174
rect -3574 222938 -3338 223174
rect -3894 222618 -3658 222854
rect -3574 222618 -3338 222854
rect -3894 186938 -3658 187174
rect -3574 186938 -3338 187174
rect -3894 186618 -3658 186854
rect -3574 186618 -3338 186854
rect -3894 150938 -3658 151174
rect -3574 150938 -3338 151174
rect -3894 150618 -3658 150854
rect -3574 150618 -3338 150854
rect -3894 114938 -3658 115174
rect -3574 114938 -3338 115174
rect -3894 114618 -3658 114854
rect -3574 114618 -3338 114854
rect -3894 78938 -3658 79174
rect -3574 78938 -3338 79174
rect -3894 78618 -3658 78854
rect -3574 78618 -3338 78854
rect -3894 42938 -3658 43174
rect -3574 42938 -3338 43174
rect -3894 42618 -3658 42854
rect -3574 42618 -3338 42854
rect -3894 6938 -3658 7174
rect -3574 6938 -3338 7174
rect -3894 6618 -3658 6854
rect -3574 6618 -3338 6854
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 669218 -2698 669454
rect -2614 669218 -2378 669454
rect -2934 668898 -2698 669134
rect -2614 668898 -2378 669134
rect -2934 633218 -2698 633454
rect -2614 633218 -2378 633454
rect -2934 632898 -2698 633134
rect -2614 632898 -2378 633134
rect -2934 597218 -2698 597454
rect -2614 597218 -2378 597454
rect -2934 596898 -2698 597134
rect -2614 596898 -2378 597134
rect -2934 561218 -2698 561454
rect -2614 561218 -2378 561454
rect -2934 560898 -2698 561134
rect -2614 560898 -2378 561134
rect -2934 525218 -2698 525454
rect -2614 525218 -2378 525454
rect -2934 524898 -2698 525134
rect -2614 524898 -2378 525134
rect -2934 489218 -2698 489454
rect -2614 489218 -2378 489454
rect -2934 488898 -2698 489134
rect -2614 488898 -2378 489134
rect -2934 453218 -2698 453454
rect -2614 453218 -2378 453454
rect -2934 452898 -2698 453134
rect -2614 452898 -2378 453134
rect -2934 417218 -2698 417454
rect -2614 417218 -2378 417454
rect -2934 416898 -2698 417134
rect -2614 416898 -2378 417134
rect -2934 381218 -2698 381454
rect -2614 381218 -2378 381454
rect -2934 380898 -2698 381134
rect -2614 380898 -2378 381134
rect -2934 345218 -2698 345454
rect -2614 345218 -2378 345454
rect -2934 344898 -2698 345134
rect -2614 344898 -2378 345134
rect -2934 309218 -2698 309454
rect -2614 309218 -2378 309454
rect -2934 308898 -2698 309134
rect -2614 308898 -2378 309134
rect -2934 273218 -2698 273454
rect -2614 273218 -2378 273454
rect -2934 272898 -2698 273134
rect -2614 272898 -2378 273134
rect -2934 237218 -2698 237454
rect -2614 237218 -2378 237454
rect -2934 236898 -2698 237134
rect -2614 236898 -2378 237134
rect -2934 201218 -2698 201454
rect -2614 201218 -2378 201454
rect -2934 200898 -2698 201134
rect -2614 200898 -2378 201134
rect -2934 165218 -2698 165454
rect -2614 165218 -2378 165454
rect -2934 164898 -2698 165134
rect -2614 164898 -2378 165134
rect -2934 129218 -2698 129454
rect -2614 129218 -2378 129454
rect -2934 128898 -2698 129134
rect -2614 128898 -2378 129134
rect -2934 93218 -2698 93454
rect -2614 93218 -2378 93454
rect -2934 92898 -2698 93134
rect -2614 92898 -2378 93134
rect -2934 57218 -2698 57454
rect -2614 57218 -2378 57454
rect -2934 56898 -2698 57134
rect -2614 56898 -2378 57134
rect -2934 21218 -2698 21454
rect -2614 21218 -2378 21454
rect -2934 20898 -2698 21134
rect -2614 20898 -2378 21134
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect 5546 -2502 5782 -2266
rect 5866 -2502 6102 -2266
rect 5546 -2822 5782 -2586
rect 5866 -2822 6102 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 9266 658658 9502 658894
rect 9586 658658 9822 658894
rect 9266 658338 9502 658574
rect 9586 658338 9822 658574
rect 9266 622658 9502 622894
rect 9586 622658 9822 622894
rect 9266 622338 9502 622574
rect 9586 622338 9822 622574
rect 9266 586658 9502 586894
rect 9586 586658 9822 586894
rect 9266 586338 9502 586574
rect 9586 586338 9822 586574
rect 9266 550658 9502 550894
rect 9586 550658 9822 550894
rect 9266 550338 9502 550574
rect 9586 550338 9822 550574
rect 9266 514658 9502 514894
rect 9586 514658 9822 514894
rect 9266 514338 9502 514574
rect 9586 514338 9822 514574
rect 9266 478658 9502 478894
rect 9586 478658 9822 478894
rect 9266 478338 9502 478574
rect 9586 478338 9822 478574
rect 9266 442658 9502 442894
rect 9586 442658 9822 442894
rect 9266 442338 9502 442574
rect 9586 442338 9822 442574
rect 9266 406658 9502 406894
rect 9586 406658 9822 406894
rect 9266 406338 9502 406574
rect 9586 406338 9822 406574
rect 9266 370658 9502 370894
rect 9586 370658 9822 370894
rect 9266 370338 9502 370574
rect 9586 370338 9822 370574
rect 9266 334658 9502 334894
rect 9586 334658 9822 334894
rect 9266 334338 9502 334574
rect 9586 334338 9822 334574
rect 9266 298658 9502 298894
rect 9586 298658 9822 298894
rect 9266 298338 9502 298574
rect 9586 298338 9822 298574
rect 9266 262658 9502 262894
rect 9586 262658 9822 262894
rect 9266 262338 9502 262574
rect 9586 262338 9822 262574
rect 9266 226658 9502 226894
rect 9586 226658 9822 226894
rect 9266 226338 9502 226574
rect 9586 226338 9822 226574
rect 9266 190658 9502 190894
rect 9586 190658 9822 190894
rect 9266 190338 9502 190574
rect 9586 190338 9822 190574
rect 9266 154658 9502 154894
rect 9586 154658 9822 154894
rect 9266 154338 9502 154574
rect 9586 154338 9822 154574
rect 9266 118658 9502 118894
rect 9586 118658 9822 118894
rect 9266 118338 9502 118574
rect 9586 118338 9822 118574
rect 9266 82658 9502 82894
rect 9586 82658 9822 82894
rect 9266 82338 9502 82574
rect 9586 82338 9822 82574
rect 9266 46658 9502 46894
rect 9586 46658 9822 46894
rect 9266 46338 9502 46574
rect 9586 46338 9822 46574
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect 9266 -4422 9502 -4186
rect 9586 -4422 9822 -4186
rect 9266 -4742 9502 -4506
rect 9586 -4742 9822 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect 30986 711322 31222 711558
rect 31306 711322 31542 711558
rect 30986 711002 31222 711238
rect 31306 711002 31542 711238
rect 27266 709402 27502 709638
rect 27586 709402 27822 709638
rect 27266 709082 27502 709318
rect 27586 709082 27822 709318
rect 23546 707482 23782 707718
rect 23866 707482 24102 707718
rect 23546 707162 23782 707398
rect 23866 707162 24102 707398
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 12986 662378 13222 662614
rect 13306 662378 13542 662614
rect 12986 662058 13222 662294
rect 13306 662058 13542 662294
rect 12986 626378 13222 626614
rect 13306 626378 13542 626614
rect 12986 626058 13222 626294
rect 13306 626058 13542 626294
rect 12986 590378 13222 590614
rect 13306 590378 13542 590614
rect 12986 590058 13222 590294
rect 13306 590058 13542 590294
rect 12986 554378 13222 554614
rect 13306 554378 13542 554614
rect 12986 554058 13222 554294
rect 13306 554058 13542 554294
rect 12986 518378 13222 518614
rect 13306 518378 13542 518614
rect 12986 518058 13222 518294
rect 13306 518058 13542 518294
rect 12986 482378 13222 482614
rect 13306 482378 13542 482614
rect 12986 482058 13222 482294
rect 13306 482058 13542 482294
rect 12986 446378 13222 446614
rect 13306 446378 13542 446614
rect 12986 446058 13222 446294
rect 13306 446058 13542 446294
rect 12986 410378 13222 410614
rect 13306 410378 13542 410614
rect 12986 410058 13222 410294
rect 13306 410058 13542 410294
rect 12986 374378 13222 374614
rect 13306 374378 13542 374614
rect 12986 374058 13222 374294
rect 13306 374058 13542 374294
rect 12986 338378 13222 338614
rect 13306 338378 13542 338614
rect 12986 338058 13222 338294
rect 13306 338058 13542 338294
rect 12986 302378 13222 302614
rect 13306 302378 13542 302614
rect 12986 302058 13222 302294
rect 13306 302058 13542 302294
rect 12986 266378 13222 266614
rect 13306 266378 13542 266614
rect 12986 266058 13222 266294
rect 13306 266058 13542 266294
rect 12986 230378 13222 230614
rect 13306 230378 13542 230614
rect 12986 230058 13222 230294
rect 13306 230058 13542 230294
rect 12986 194378 13222 194614
rect 13306 194378 13542 194614
rect 12986 194058 13222 194294
rect 13306 194058 13542 194294
rect 12986 158378 13222 158614
rect 13306 158378 13542 158614
rect 12986 158058 13222 158294
rect 13306 158058 13542 158294
rect 12986 122378 13222 122614
rect 13306 122378 13542 122614
rect 12986 122058 13222 122294
rect 13306 122058 13542 122294
rect 12986 86378 13222 86614
rect 13306 86378 13542 86614
rect 12986 86058 13222 86294
rect 13306 86058 13542 86294
rect 12986 50378 13222 50614
rect 13306 50378 13542 50614
rect 12986 50058 13222 50294
rect 13306 50058 13542 50294
rect 12986 14378 13222 14614
rect 13306 14378 13542 14614
rect 12986 14058 13222 14294
rect 13306 14058 13542 14294
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect 19826 705562 20062 705798
rect 20146 705562 20382 705798
rect 19826 705242 20062 705478
rect 20146 705242 20382 705478
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -1542 20062 -1306
rect 20146 -1542 20382 -1306
rect 19826 -1862 20062 -1626
rect 20146 -1862 20382 -1626
rect 23546 672938 23782 673174
rect 23866 672938 24102 673174
rect 23546 672618 23782 672854
rect 23866 672618 24102 672854
rect 23546 636938 23782 637174
rect 23866 636938 24102 637174
rect 23546 636618 23782 636854
rect 23866 636618 24102 636854
rect 23546 600938 23782 601174
rect 23866 600938 24102 601174
rect 23546 600618 23782 600854
rect 23866 600618 24102 600854
rect 23546 564938 23782 565174
rect 23866 564938 24102 565174
rect 23546 564618 23782 564854
rect 23866 564618 24102 564854
rect 23546 528938 23782 529174
rect 23866 528938 24102 529174
rect 23546 528618 23782 528854
rect 23866 528618 24102 528854
rect 23546 492938 23782 493174
rect 23866 492938 24102 493174
rect 23546 492618 23782 492854
rect 23866 492618 24102 492854
rect 23546 456938 23782 457174
rect 23866 456938 24102 457174
rect 23546 456618 23782 456854
rect 23866 456618 24102 456854
rect 23546 420938 23782 421174
rect 23866 420938 24102 421174
rect 23546 420618 23782 420854
rect 23866 420618 24102 420854
rect 23546 384938 23782 385174
rect 23866 384938 24102 385174
rect 23546 384618 23782 384854
rect 23866 384618 24102 384854
rect 23546 348938 23782 349174
rect 23866 348938 24102 349174
rect 23546 348618 23782 348854
rect 23866 348618 24102 348854
rect 23546 312938 23782 313174
rect 23866 312938 24102 313174
rect 23546 312618 23782 312854
rect 23866 312618 24102 312854
rect 23546 276938 23782 277174
rect 23866 276938 24102 277174
rect 23546 276618 23782 276854
rect 23866 276618 24102 276854
rect 23546 240938 23782 241174
rect 23866 240938 24102 241174
rect 23546 240618 23782 240854
rect 23866 240618 24102 240854
rect 23546 204938 23782 205174
rect 23866 204938 24102 205174
rect 23546 204618 23782 204854
rect 23866 204618 24102 204854
rect 23546 168938 23782 169174
rect 23866 168938 24102 169174
rect 23546 168618 23782 168854
rect 23866 168618 24102 168854
rect 23546 132938 23782 133174
rect 23866 132938 24102 133174
rect 23546 132618 23782 132854
rect 23866 132618 24102 132854
rect 23546 96938 23782 97174
rect 23866 96938 24102 97174
rect 23546 96618 23782 96854
rect 23866 96618 24102 96854
rect 23546 60938 23782 61174
rect 23866 60938 24102 61174
rect 23546 60618 23782 60854
rect 23866 60618 24102 60854
rect 23546 24938 23782 25174
rect 23866 24938 24102 25174
rect 23546 24618 23782 24854
rect 23866 24618 24102 24854
rect 23546 -3462 23782 -3226
rect 23866 -3462 24102 -3226
rect 23546 -3782 23782 -3546
rect 23866 -3782 24102 -3546
rect 27266 676658 27502 676894
rect 27586 676658 27822 676894
rect 27266 676338 27502 676574
rect 27586 676338 27822 676574
rect 27266 640658 27502 640894
rect 27586 640658 27822 640894
rect 27266 640338 27502 640574
rect 27586 640338 27822 640574
rect 27266 604658 27502 604894
rect 27586 604658 27822 604894
rect 27266 604338 27502 604574
rect 27586 604338 27822 604574
rect 27266 568658 27502 568894
rect 27586 568658 27822 568894
rect 27266 568338 27502 568574
rect 27586 568338 27822 568574
rect 27266 532658 27502 532894
rect 27586 532658 27822 532894
rect 27266 532338 27502 532574
rect 27586 532338 27822 532574
rect 27266 496658 27502 496894
rect 27586 496658 27822 496894
rect 27266 496338 27502 496574
rect 27586 496338 27822 496574
rect 27266 460658 27502 460894
rect 27586 460658 27822 460894
rect 27266 460338 27502 460574
rect 27586 460338 27822 460574
rect 27266 424658 27502 424894
rect 27586 424658 27822 424894
rect 27266 424338 27502 424574
rect 27586 424338 27822 424574
rect 27266 388658 27502 388894
rect 27586 388658 27822 388894
rect 27266 388338 27502 388574
rect 27586 388338 27822 388574
rect 27266 352658 27502 352894
rect 27586 352658 27822 352894
rect 27266 352338 27502 352574
rect 27586 352338 27822 352574
rect 27266 316658 27502 316894
rect 27586 316658 27822 316894
rect 27266 316338 27502 316574
rect 27586 316338 27822 316574
rect 27266 280658 27502 280894
rect 27586 280658 27822 280894
rect 27266 280338 27502 280574
rect 27586 280338 27822 280574
rect 27266 244658 27502 244894
rect 27586 244658 27822 244894
rect 27266 244338 27502 244574
rect 27586 244338 27822 244574
rect 27266 208658 27502 208894
rect 27586 208658 27822 208894
rect 27266 208338 27502 208574
rect 27586 208338 27822 208574
rect 27266 172658 27502 172894
rect 27586 172658 27822 172894
rect 27266 172338 27502 172574
rect 27586 172338 27822 172574
rect 27266 136658 27502 136894
rect 27586 136658 27822 136894
rect 27266 136338 27502 136574
rect 27586 136338 27822 136574
rect 27266 100658 27502 100894
rect 27586 100658 27822 100894
rect 27266 100338 27502 100574
rect 27586 100338 27822 100574
rect 27266 64658 27502 64894
rect 27586 64658 27822 64894
rect 27266 64338 27502 64574
rect 27586 64338 27822 64574
rect 27266 28658 27502 28894
rect 27586 28658 27822 28894
rect 27266 28338 27502 28574
rect 27586 28338 27822 28574
rect 27266 -5382 27502 -5146
rect 27586 -5382 27822 -5146
rect 27266 -5702 27502 -5466
rect 27586 -5702 27822 -5466
rect 48986 710362 49222 710598
rect 49306 710362 49542 710598
rect 48986 710042 49222 710278
rect 49306 710042 49542 710278
rect 45266 708442 45502 708678
rect 45586 708442 45822 708678
rect 45266 708122 45502 708358
rect 45586 708122 45822 708358
rect 41546 706522 41782 706758
rect 41866 706522 42102 706758
rect 41546 706202 41782 706438
rect 41866 706202 42102 706438
rect 30986 680378 31222 680614
rect 31306 680378 31542 680614
rect 30986 680058 31222 680294
rect 31306 680058 31542 680294
rect 30986 644378 31222 644614
rect 31306 644378 31542 644614
rect 30986 644058 31222 644294
rect 31306 644058 31542 644294
rect 30986 608378 31222 608614
rect 31306 608378 31542 608614
rect 30986 608058 31222 608294
rect 31306 608058 31542 608294
rect 30986 572378 31222 572614
rect 31306 572378 31542 572614
rect 30986 572058 31222 572294
rect 31306 572058 31542 572294
rect 30986 536378 31222 536614
rect 31306 536378 31542 536614
rect 30986 536058 31222 536294
rect 31306 536058 31542 536294
rect 30986 500378 31222 500614
rect 31306 500378 31542 500614
rect 30986 500058 31222 500294
rect 31306 500058 31542 500294
rect 30986 464378 31222 464614
rect 31306 464378 31542 464614
rect 30986 464058 31222 464294
rect 31306 464058 31542 464294
rect 30986 428378 31222 428614
rect 31306 428378 31542 428614
rect 30986 428058 31222 428294
rect 31306 428058 31542 428294
rect 30986 392378 31222 392614
rect 31306 392378 31542 392614
rect 30986 392058 31222 392294
rect 31306 392058 31542 392294
rect 30986 356378 31222 356614
rect 31306 356378 31542 356614
rect 30986 356058 31222 356294
rect 31306 356058 31542 356294
rect 30986 320378 31222 320614
rect 31306 320378 31542 320614
rect 30986 320058 31222 320294
rect 31306 320058 31542 320294
rect 30986 284378 31222 284614
rect 31306 284378 31542 284614
rect 30986 284058 31222 284294
rect 31306 284058 31542 284294
rect 30986 248378 31222 248614
rect 31306 248378 31542 248614
rect 30986 248058 31222 248294
rect 31306 248058 31542 248294
rect 30986 212378 31222 212614
rect 31306 212378 31542 212614
rect 30986 212058 31222 212294
rect 31306 212058 31542 212294
rect 30986 176378 31222 176614
rect 31306 176378 31542 176614
rect 30986 176058 31222 176294
rect 31306 176058 31542 176294
rect 30986 140378 31222 140614
rect 31306 140378 31542 140614
rect 30986 140058 31222 140294
rect 31306 140058 31542 140294
rect 30986 104378 31222 104614
rect 31306 104378 31542 104614
rect 30986 104058 31222 104294
rect 31306 104058 31542 104294
rect 30986 68378 31222 68614
rect 31306 68378 31542 68614
rect 30986 68058 31222 68294
rect 31306 68058 31542 68294
rect 30986 32378 31222 32614
rect 31306 32378 31542 32614
rect 30986 32058 31222 32294
rect 31306 32058 31542 32294
rect 12986 -6342 13222 -6106
rect 13306 -6342 13542 -6106
rect 12986 -6662 13222 -6426
rect 13306 -6662 13542 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 41546 654938 41782 655174
rect 41866 654938 42102 655174
rect 41546 654618 41782 654854
rect 41866 654618 42102 654854
rect 41546 618938 41782 619174
rect 41866 618938 42102 619174
rect 41546 618618 41782 618854
rect 41866 618618 42102 618854
rect 41546 582938 41782 583174
rect 41866 582938 42102 583174
rect 41546 582618 41782 582854
rect 41866 582618 42102 582854
rect 41546 546938 41782 547174
rect 41866 546938 42102 547174
rect 41546 546618 41782 546854
rect 41866 546618 42102 546854
rect 41546 510938 41782 511174
rect 41866 510938 42102 511174
rect 41546 510618 41782 510854
rect 41866 510618 42102 510854
rect 41546 474938 41782 475174
rect 41866 474938 42102 475174
rect 41546 474618 41782 474854
rect 41866 474618 42102 474854
rect 41546 438938 41782 439174
rect 41866 438938 42102 439174
rect 41546 438618 41782 438854
rect 41866 438618 42102 438854
rect 41546 402938 41782 403174
rect 41866 402938 42102 403174
rect 41546 402618 41782 402854
rect 41866 402618 42102 402854
rect 41546 366938 41782 367174
rect 41866 366938 42102 367174
rect 41546 366618 41782 366854
rect 41866 366618 42102 366854
rect 41546 330938 41782 331174
rect 41866 330938 42102 331174
rect 41546 330618 41782 330854
rect 41866 330618 42102 330854
rect 41546 294938 41782 295174
rect 41866 294938 42102 295174
rect 41546 294618 41782 294854
rect 41866 294618 42102 294854
rect 41546 258938 41782 259174
rect 41866 258938 42102 259174
rect 41546 258618 41782 258854
rect 41866 258618 42102 258854
rect 41546 222938 41782 223174
rect 41866 222938 42102 223174
rect 41546 222618 41782 222854
rect 41866 222618 42102 222854
rect 41546 186938 41782 187174
rect 41866 186938 42102 187174
rect 41546 186618 41782 186854
rect 41866 186618 42102 186854
rect 41546 150938 41782 151174
rect 41866 150938 42102 151174
rect 41546 150618 41782 150854
rect 41866 150618 42102 150854
rect 41546 114938 41782 115174
rect 41866 114938 42102 115174
rect 41546 114618 41782 114854
rect 41866 114618 42102 114854
rect 41546 78938 41782 79174
rect 41866 78938 42102 79174
rect 41546 78618 41782 78854
rect 41866 78618 42102 78854
rect 41546 42938 41782 43174
rect 41866 42938 42102 43174
rect 41546 42618 41782 42854
rect 41866 42618 42102 42854
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -2502 41782 -2266
rect 41866 -2502 42102 -2266
rect 41546 -2822 41782 -2586
rect 41866 -2822 42102 -2586
rect 45266 694658 45502 694894
rect 45586 694658 45822 694894
rect 45266 694338 45502 694574
rect 45586 694338 45822 694574
rect 45266 658658 45502 658894
rect 45586 658658 45822 658894
rect 45266 658338 45502 658574
rect 45586 658338 45822 658574
rect 45266 622658 45502 622894
rect 45586 622658 45822 622894
rect 45266 622338 45502 622574
rect 45586 622338 45822 622574
rect 45266 586658 45502 586894
rect 45586 586658 45822 586894
rect 45266 586338 45502 586574
rect 45586 586338 45822 586574
rect 45266 550658 45502 550894
rect 45586 550658 45822 550894
rect 45266 550338 45502 550574
rect 45586 550338 45822 550574
rect 45266 514658 45502 514894
rect 45586 514658 45822 514894
rect 45266 514338 45502 514574
rect 45586 514338 45822 514574
rect 45266 478658 45502 478894
rect 45586 478658 45822 478894
rect 45266 478338 45502 478574
rect 45586 478338 45822 478574
rect 66986 711322 67222 711558
rect 67306 711322 67542 711558
rect 66986 711002 67222 711238
rect 67306 711002 67542 711238
rect 63266 709402 63502 709638
rect 63586 709402 63822 709638
rect 63266 709082 63502 709318
rect 63586 709082 63822 709318
rect 59546 707482 59782 707718
rect 59866 707482 60102 707718
rect 59546 707162 59782 707398
rect 59866 707162 60102 707398
rect 48986 698378 49222 698614
rect 49306 698378 49542 698614
rect 48986 698058 49222 698294
rect 49306 698058 49542 698294
rect 48986 662378 49222 662614
rect 49306 662378 49542 662614
rect 48986 662058 49222 662294
rect 49306 662058 49542 662294
rect 48986 626378 49222 626614
rect 49306 626378 49542 626614
rect 48986 626058 49222 626294
rect 49306 626058 49542 626294
rect 48986 590378 49222 590614
rect 49306 590378 49542 590614
rect 48986 590058 49222 590294
rect 49306 590058 49542 590294
rect 48986 554378 49222 554614
rect 49306 554378 49542 554614
rect 48986 554058 49222 554294
rect 49306 554058 49542 554294
rect 48986 518378 49222 518614
rect 49306 518378 49542 518614
rect 48986 518058 49222 518294
rect 49306 518058 49542 518294
rect 48986 482378 49222 482614
rect 49306 482378 49542 482614
rect 48986 482058 49222 482294
rect 49306 482058 49542 482294
rect 55826 705562 56062 705798
rect 56146 705562 56382 705798
rect 55826 705242 56062 705478
rect 56146 705242 56382 705478
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 59546 672938 59782 673174
rect 59866 672938 60102 673174
rect 59546 672618 59782 672854
rect 59866 672618 60102 672854
rect 59546 636938 59782 637174
rect 59866 636938 60102 637174
rect 59546 636618 59782 636854
rect 59866 636618 60102 636854
rect 59546 600938 59782 601174
rect 59866 600938 60102 601174
rect 59546 600618 59782 600854
rect 59866 600618 60102 600854
rect 59546 564938 59782 565174
rect 59866 564938 60102 565174
rect 59546 564618 59782 564854
rect 59866 564618 60102 564854
rect 59546 528938 59782 529174
rect 59866 528938 60102 529174
rect 59546 528618 59782 528854
rect 59866 528618 60102 528854
rect 59546 492938 59782 493174
rect 59866 492938 60102 493174
rect 59546 492618 59782 492854
rect 59866 492618 60102 492854
rect 63266 676658 63502 676894
rect 63586 676658 63822 676894
rect 63266 676338 63502 676574
rect 63586 676338 63822 676574
rect 63266 640658 63502 640894
rect 63586 640658 63822 640894
rect 63266 640338 63502 640574
rect 63586 640338 63822 640574
rect 63266 604658 63502 604894
rect 63586 604658 63822 604894
rect 63266 604338 63502 604574
rect 63586 604338 63822 604574
rect 63266 568658 63502 568894
rect 63586 568658 63822 568894
rect 63266 568338 63502 568574
rect 63586 568338 63822 568574
rect 63266 532658 63502 532894
rect 63586 532658 63822 532894
rect 63266 532338 63502 532574
rect 63586 532338 63822 532574
rect 63266 496658 63502 496894
rect 63586 496658 63822 496894
rect 63266 496338 63502 496574
rect 63586 496338 63822 496574
rect 84986 710362 85222 710598
rect 85306 710362 85542 710598
rect 84986 710042 85222 710278
rect 85306 710042 85542 710278
rect 81266 708442 81502 708678
rect 81586 708442 81822 708678
rect 81266 708122 81502 708358
rect 81586 708122 81822 708358
rect 77546 706522 77782 706758
rect 77866 706522 78102 706758
rect 77546 706202 77782 706438
rect 77866 706202 78102 706438
rect 66986 680378 67222 680614
rect 67306 680378 67542 680614
rect 66986 680058 67222 680294
rect 67306 680058 67542 680294
rect 66986 644378 67222 644614
rect 67306 644378 67542 644614
rect 66986 644058 67222 644294
rect 67306 644058 67542 644294
rect 66986 608378 67222 608614
rect 67306 608378 67542 608614
rect 66986 608058 67222 608294
rect 67306 608058 67542 608294
rect 66986 572378 67222 572614
rect 67306 572378 67542 572614
rect 66986 572058 67222 572294
rect 67306 572058 67542 572294
rect 66986 536378 67222 536614
rect 67306 536378 67542 536614
rect 66986 536058 67222 536294
rect 67306 536058 67542 536294
rect 66986 500378 67222 500614
rect 67306 500378 67542 500614
rect 66986 500058 67222 500294
rect 67306 500058 67542 500294
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 73826 579218 74062 579454
rect 74146 579218 74382 579454
rect 73826 578898 74062 579134
rect 74146 578898 74382 579134
rect 73826 543218 74062 543454
rect 74146 543218 74382 543454
rect 73826 542898 74062 543134
rect 74146 542898 74382 543134
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 77546 654938 77782 655174
rect 77866 654938 78102 655174
rect 77546 654618 77782 654854
rect 77866 654618 78102 654854
rect 77546 618938 77782 619174
rect 77866 618938 78102 619174
rect 77546 618618 77782 618854
rect 77866 618618 78102 618854
rect 77546 582938 77782 583174
rect 77866 582938 78102 583174
rect 77546 582618 77782 582854
rect 77866 582618 78102 582854
rect 77546 546938 77782 547174
rect 77866 546938 78102 547174
rect 77546 546618 77782 546854
rect 77866 546618 78102 546854
rect 77546 510938 77782 511174
rect 77866 510938 78102 511174
rect 77546 510618 77782 510854
rect 77866 510618 78102 510854
rect 77546 474938 77782 475174
rect 77866 474938 78102 475174
rect 77546 474618 77782 474854
rect 77866 474618 78102 474854
rect 81266 694658 81502 694894
rect 81586 694658 81822 694894
rect 81266 694338 81502 694574
rect 81586 694338 81822 694574
rect 81266 658658 81502 658894
rect 81586 658658 81822 658894
rect 81266 658338 81502 658574
rect 81586 658338 81822 658574
rect 81266 622658 81502 622894
rect 81586 622658 81822 622894
rect 81266 622338 81502 622574
rect 81586 622338 81822 622574
rect 81266 586658 81502 586894
rect 81586 586658 81822 586894
rect 81266 586338 81502 586574
rect 81586 586338 81822 586574
rect 81266 550658 81502 550894
rect 81586 550658 81822 550894
rect 81266 550338 81502 550574
rect 81586 550338 81822 550574
rect 81266 514658 81502 514894
rect 81586 514658 81822 514894
rect 81266 514338 81502 514574
rect 81586 514338 81822 514574
rect 81266 478658 81502 478894
rect 81586 478658 81822 478894
rect 81266 478338 81502 478574
rect 81586 478338 81822 478574
rect 102986 711322 103222 711558
rect 103306 711322 103542 711558
rect 102986 711002 103222 711238
rect 103306 711002 103542 711238
rect 99266 709402 99502 709638
rect 99586 709402 99822 709638
rect 99266 709082 99502 709318
rect 99586 709082 99822 709318
rect 95546 707482 95782 707718
rect 95866 707482 96102 707718
rect 95546 707162 95782 707398
rect 95866 707162 96102 707398
rect 84986 698378 85222 698614
rect 85306 698378 85542 698614
rect 84986 698058 85222 698294
rect 85306 698058 85542 698294
rect 84986 662378 85222 662614
rect 85306 662378 85542 662614
rect 84986 662058 85222 662294
rect 85306 662058 85542 662294
rect 84986 626378 85222 626614
rect 85306 626378 85542 626614
rect 84986 626058 85222 626294
rect 85306 626058 85542 626294
rect 84986 590378 85222 590614
rect 85306 590378 85542 590614
rect 84986 590058 85222 590294
rect 85306 590058 85542 590294
rect 84986 554378 85222 554614
rect 85306 554378 85542 554614
rect 84986 554058 85222 554294
rect 85306 554058 85542 554294
rect 84986 518378 85222 518614
rect 85306 518378 85542 518614
rect 84986 518058 85222 518294
rect 85306 518058 85542 518294
rect 84986 482378 85222 482614
rect 85306 482378 85542 482614
rect 84986 482058 85222 482294
rect 85306 482058 85542 482294
rect 91826 705562 92062 705798
rect 92146 705562 92382 705798
rect 91826 705242 92062 705478
rect 92146 705242 92382 705478
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 91826 561218 92062 561454
rect 92146 561218 92382 561454
rect 91826 560898 92062 561134
rect 92146 560898 92382 561134
rect 91826 525218 92062 525454
rect 92146 525218 92382 525454
rect 91826 524898 92062 525134
rect 92146 524898 92382 525134
rect 91826 489218 92062 489454
rect 92146 489218 92382 489454
rect 91826 488898 92062 489134
rect 92146 488898 92382 489134
rect 95546 672938 95782 673174
rect 95866 672938 96102 673174
rect 95546 672618 95782 672854
rect 95866 672618 96102 672854
rect 95546 636938 95782 637174
rect 95866 636938 96102 637174
rect 95546 636618 95782 636854
rect 95866 636618 96102 636854
rect 95546 600938 95782 601174
rect 95866 600938 96102 601174
rect 95546 600618 95782 600854
rect 95866 600618 96102 600854
rect 95546 564938 95782 565174
rect 95866 564938 96102 565174
rect 95546 564618 95782 564854
rect 95866 564618 96102 564854
rect 95546 528938 95782 529174
rect 95866 528938 96102 529174
rect 95546 528618 95782 528854
rect 95866 528618 96102 528854
rect 95546 492938 95782 493174
rect 95866 492938 96102 493174
rect 95546 492618 95782 492854
rect 95866 492618 96102 492854
rect 99266 676658 99502 676894
rect 99586 676658 99822 676894
rect 99266 676338 99502 676574
rect 99586 676338 99822 676574
rect 99266 640658 99502 640894
rect 99586 640658 99822 640894
rect 99266 640338 99502 640574
rect 99586 640338 99822 640574
rect 99266 604658 99502 604894
rect 99586 604658 99822 604894
rect 99266 604338 99502 604574
rect 99586 604338 99822 604574
rect 99266 568658 99502 568894
rect 99586 568658 99822 568894
rect 99266 568338 99502 568574
rect 99586 568338 99822 568574
rect 99266 532658 99502 532894
rect 99586 532658 99822 532894
rect 99266 532338 99502 532574
rect 99586 532338 99822 532574
rect 99266 496658 99502 496894
rect 99586 496658 99822 496894
rect 99266 496338 99502 496574
rect 99586 496338 99822 496574
rect 120986 710362 121222 710598
rect 121306 710362 121542 710598
rect 120986 710042 121222 710278
rect 121306 710042 121542 710278
rect 117266 708442 117502 708678
rect 117586 708442 117822 708678
rect 117266 708122 117502 708358
rect 117586 708122 117822 708358
rect 113546 706522 113782 706758
rect 113866 706522 114102 706758
rect 113546 706202 113782 706438
rect 113866 706202 114102 706438
rect 102986 680378 103222 680614
rect 103306 680378 103542 680614
rect 102986 680058 103222 680294
rect 103306 680058 103542 680294
rect 102986 644378 103222 644614
rect 103306 644378 103542 644614
rect 102986 644058 103222 644294
rect 103306 644058 103542 644294
rect 102986 608378 103222 608614
rect 103306 608378 103542 608614
rect 102986 608058 103222 608294
rect 103306 608058 103542 608294
rect 102986 572378 103222 572614
rect 103306 572378 103542 572614
rect 102986 572058 103222 572294
rect 103306 572058 103542 572294
rect 102986 536378 103222 536614
rect 103306 536378 103542 536614
rect 102986 536058 103222 536294
rect 103306 536058 103542 536294
rect 102986 500378 103222 500614
rect 103306 500378 103542 500614
rect 102986 500058 103222 500294
rect 103306 500058 103542 500294
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 109826 507218 110062 507454
rect 110146 507218 110382 507454
rect 109826 506898 110062 507134
rect 110146 506898 110382 507134
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 113546 654938 113782 655174
rect 113866 654938 114102 655174
rect 113546 654618 113782 654854
rect 113866 654618 114102 654854
rect 113546 618938 113782 619174
rect 113866 618938 114102 619174
rect 113546 618618 113782 618854
rect 113866 618618 114102 618854
rect 113546 582938 113782 583174
rect 113866 582938 114102 583174
rect 113546 582618 113782 582854
rect 113866 582618 114102 582854
rect 113546 546938 113782 547174
rect 113866 546938 114102 547174
rect 113546 546618 113782 546854
rect 113866 546618 114102 546854
rect 113546 510938 113782 511174
rect 113866 510938 114102 511174
rect 113546 510618 113782 510854
rect 113866 510618 114102 510854
rect 113546 474938 113782 475174
rect 113866 474938 114102 475174
rect 113546 474618 113782 474854
rect 113866 474618 114102 474854
rect 117266 694658 117502 694894
rect 117586 694658 117822 694894
rect 117266 694338 117502 694574
rect 117586 694338 117822 694574
rect 117266 658658 117502 658894
rect 117586 658658 117822 658894
rect 117266 658338 117502 658574
rect 117586 658338 117822 658574
rect 117266 622658 117502 622894
rect 117586 622658 117822 622894
rect 117266 622338 117502 622574
rect 117586 622338 117822 622574
rect 117266 586658 117502 586894
rect 117586 586658 117822 586894
rect 117266 586338 117502 586574
rect 117586 586338 117822 586574
rect 117266 550658 117502 550894
rect 117586 550658 117822 550894
rect 117266 550338 117502 550574
rect 117586 550338 117822 550574
rect 117266 514658 117502 514894
rect 117586 514658 117822 514894
rect 117266 514338 117502 514574
rect 117586 514338 117822 514574
rect 117266 478658 117502 478894
rect 117586 478658 117822 478894
rect 117266 478338 117502 478574
rect 117586 478338 117822 478574
rect 138986 711322 139222 711558
rect 139306 711322 139542 711558
rect 138986 711002 139222 711238
rect 139306 711002 139542 711238
rect 135266 709402 135502 709638
rect 135586 709402 135822 709638
rect 135266 709082 135502 709318
rect 135586 709082 135822 709318
rect 131546 707482 131782 707718
rect 131866 707482 132102 707718
rect 131546 707162 131782 707398
rect 131866 707162 132102 707398
rect 120986 698378 121222 698614
rect 121306 698378 121542 698614
rect 120986 698058 121222 698294
rect 121306 698058 121542 698294
rect 120986 662378 121222 662614
rect 121306 662378 121542 662614
rect 120986 662058 121222 662294
rect 121306 662058 121542 662294
rect 120986 626378 121222 626614
rect 121306 626378 121542 626614
rect 120986 626058 121222 626294
rect 121306 626058 121542 626294
rect 120986 590378 121222 590614
rect 121306 590378 121542 590614
rect 120986 590058 121222 590294
rect 121306 590058 121542 590294
rect 120986 554378 121222 554614
rect 121306 554378 121542 554614
rect 120986 554058 121222 554294
rect 121306 554058 121542 554294
rect 120986 518378 121222 518614
rect 121306 518378 121542 518614
rect 120986 518058 121222 518294
rect 121306 518058 121542 518294
rect 120986 482378 121222 482614
rect 121306 482378 121542 482614
rect 120986 482058 121222 482294
rect 121306 482058 121542 482294
rect 127826 705562 128062 705798
rect 128146 705562 128382 705798
rect 127826 705242 128062 705478
rect 128146 705242 128382 705478
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 127826 525218 128062 525454
rect 128146 525218 128382 525454
rect 127826 524898 128062 525134
rect 128146 524898 128382 525134
rect 127826 489218 128062 489454
rect 128146 489218 128382 489454
rect 127826 488898 128062 489134
rect 128146 488898 128382 489134
rect 131546 672938 131782 673174
rect 131866 672938 132102 673174
rect 131546 672618 131782 672854
rect 131866 672618 132102 672854
rect 131546 636938 131782 637174
rect 131866 636938 132102 637174
rect 131546 636618 131782 636854
rect 131866 636618 132102 636854
rect 131546 600938 131782 601174
rect 131866 600938 132102 601174
rect 131546 600618 131782 600854
rect 131866 600618 132102 600854
rect 131546 564938 131782 565174
rect 131866 564938 132102 565174
rect 131546 564618 131782 564854
rect 131866 564618 132102 564854
rect 131546 528938 131782 529174
rect 131866 528938 132102 529174
rect 131546 528618 131782 528854
rect 131866 528618 132102 528854
rect 131546 492938 131782 493174
rect 131866 492938 132102 493174
rect 131546 492618 131782 492854
rect 131866 492618 132102 492854
rect 135266 676658 135502 676894
rect 135586 676658 135822 676894
rect 135266 676338 135502 676574
rect 135586 676338 135822 676574
rect 135266 640658 135502 640894
rect 135586 640658 135822 640894
rect 135266 640338 135502 640574
rect 135586 640338 135822 640574
rect 135266 604658 135502 604894
rect 135586 604658 135822 604894
rect 135266 604338 135502 604574
rect 135586 604338 135822 604574
rect 135266 568658 135502 568894
rect 135586 568658 135822 568894
rect 135266 568338 135502 568574
rect 135586 568338 135822 568574
rect 135266 532658 135502 532894
rect 135586 532658 135822 532894
rect 135266 532338 135502 532574
rect 135586 532338 135822 532574
rect 135266 496658 135502 496894
rect 135586 496658 135822 496894
rect 135266 496338 135502 496574
rect 135586 496338 135822 496574
rect 156986 710362 157222 710598
rect 157306 710362 157542 710598
rect 156986 710042 157222 710278
rect 157306 710042 157542 710278
rect 153266 708442 153502 708678
rect 153586 708442 153822 708678
rect 153266 708122 153502 708358
rect 153586 708122 153822 708358
rect 149546 706522 149782 706758
rect 149866 706522 150102 706758
rect 149546 706202 149782 706438
rect 149866 706202 150102 706438
rect 138986 680378 139222 680614
rect 139306 680378 139542 680614
rect 138986 680058 139222 680294
rect 139306 680058 139542 680294
rect 138986 644378 139222 644614
rect 139306 644378 139542 644614
rect 138986 644058 139222 644294
rect 139306 644058 139542 644294
rect 138986 608378 139222 608614
rect 139306 608378 139542 608614
rect 138986 608058 139222 608294
rect 139306 608058 139542 608294
rect 138986 572378 139222 572614
rect 139306 572378 139542 572614
rect 138986 572058 139222 572294
rect 139306 572058 139542 572294
rect 138986 536378 139222 536614
rect 139306 536378 139542 536614
rect 138986 536058 139222 536294
rect 139306 536058 139542 536294
rect 138986 500378 139222 500614
rect 139306 500378 139542 500614
rect 138986 500058 139222 500294
rect 139306 500058 139542 500294
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 149546 654938 149782 655174
rect 149866 654938 150102 655174
rect 149546 654618 149782 654854
rect 149866 654618 150102 654854
rect 149546 618938 149782 619174
rect 149866 618938 150102 619174
rect 149546 618618 149782 618854
rect 149866 618618 150102 618854
rect 149546 582938 149782 583174
rect 149866 582938 150102 583174
rect 149546 582618 149782 582854
rect 149866 582618 150102 582854
rect 149546 546938 149782 547174
rect 149866 546938 150102 547174
rect 149546 546618 149782 546854
rect 149866 546618 150102 546854
rect 149546 510938 149782 511174
rect 149866 510938 150102 511174
rect 149546 510618 149782 510854
rect 149866 510618 150102 510854
rect 149546 474938 149782 475174
rect 149866 474938 150102 475174
rect 149546 474618 149782 474854
rect 149866 474618 150102 474854
rect 153266 694658 153502 694894
rect 153586 694658 153822 694894
rect 153266 694338 153502 694574
rect 153586 694338 153822 694574
rect 153266 658658 153502 658894
rect 153586 658658 153822 658894
rect 153266 658338 153502 658574
rect 153586 658338 153822 658574
rect 153266 622658 153502 622894
rect 153586 622658 153822 622894
rect 153266 622338 153502 622574
rect 153586 622338 153822 622574
rect 153266 586658 153502 586894
rect 153586 586658 153822 586894
rect 153266 586338 153502 586574
rect 153586 586338 153822 586574
rect 153266 550658 153502 550894
rect 153586 550658 153822 550894
rect 153266 550338 153502 550574
rect 153586 550338 153822 550574
rect 153266 514658 153502 514894
rect 153586 514658 153822 514894
rect 153266 514338 153502 514574
rect 153586 514338 153822 514574
rect 153266 478658 153502 478894
rect 153586 478658 153822 478894
rect 153266 478338 153502 478574
rect 153586 478338 153822 478574
rect 174986 711322 175222 711558
rect 175306 711322 175542 711558
rect 174986 711002 175222 711238
rect 175306 711002 175542 711238
rect 171266 709402 171502 709638
rect 171586 709402 171822 709638
rect 171266 709082 171502 709318
rect 171586 709082 171822 709318
rect 167546 707482 167782 707718
rect 167866 707482 168102 707718
rect 167546 707162 167782 707398
rect 167866 707162 168102 707398
rect 156986 698378 157222 698614
rect 157306 698378 157542 698614
rect 156986 698058 157222 698294
rect 157306 698058 157542 698294
rect 156986 662378 157222 662614
rect 157306 662378 157542 662614
rect 156986 662058 157222 662294
rect 157306 662058 157542 662294
rect 156986 626378 157222 626614
rect 157306 626378 157542 626614
rect 156986 626058 157222 626294
rect 157306 626058 157542 626294
rect 156986 590378 157222 590614
rect 157306 590378 157542 590614
rect 156986 590058 157222 590294
rect 157306 590058 157542 590294
rect 156986 554378 157222 554614
rect 157306 554378 157542 554614
rect 156986 554058 157222 554294
rect 157306 554058 157542 554294
rect 156986 518378 157222 518614
rect 157306 518378 157542 518614
rect 156986 518058 157222 518294
rect 157306 518058 157542 518294
rect 156986 482378 157222 482614
rect 157306 482378 157542 482614
rect 156986 482058 157222 482294
rect 157306 482058 157542 482294
rect 163826 705562 164062 705798
rect 164146 705562 164382 705798
rect 163826 705242 164062 705478
rect 164146 705242 164382 705478
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 163826 561218 164062 561454
rect 164146 561218 164382 561454
rect 163826 560898 164062 561134
rect 164146 560898 164382 561134
rect 163826 525218 164062 525454
rect 164146 525218 164382 525454
rect 163826 524898 164062 525134
rect 164146 524898 164382 525134
rect 163826 489218 164062 489454
rect 164146 489218 164382 489454
rect 163826 488898 164062 489134
rect 164146 488898 164382 489134
rect 167546 672938 167782 673174
rect 167866 672938 168102 673174
rect 167546 672618 167782 672854
rect 167866 672618 168102 672854
rect 167546 636938 167782 637174
rect 167866 636938 168102 637174
rect 167546 636618 167782 636854
rect 167866 636618 168102 636854
rect 167546 600938 167782 601174
rect 167866 600938 168102 601174
rect 167546 600618 167782 600854
rect 167866 600618 168102 600854
rect 167546 564938 167782 565174
rect 167866 564938 168102 565174
rect 167546 564618 167782 564854
rect 167866 564618 168102 564854
rect 167546 528938 167782 529174
rect 167866 528938 168102 529174
rect 167546 528618 167782 528854
rect 167866 528618 168102 528854
rect 167546 492938 167782 493174
rect 167866 492938 168102 493174
rect 167546 492618 167782 492854
rect 167866 492618 168102 492854
rect 171266 676658 171502 676894
rect 171586 676658 171822 676894
rect 171266 676338 171502 676574
rect 171586 676338 171822 676574
rect 171266 640658 171502 640894
rect 171586 640658 171822 640894
rect 171266 640338 171502 640574
rect 171586 640338 171822 640574
rect 171266 604658 171502 604894
rect 171586 604658 171822 604894
rect 171266 604338 171502 604574
rect 171586 604338 171822 604574
rect 171266 568658 171502 568894
rect 171586 568658 171822 568894
rect 171266 568338 171502 568574
rect 171586 568338 171822 568574
rect 171266 532658 171502 532894
rect 171586 532658 171822 532894
rect 171266 532338 171502 532574
rect 171586 532338 171822 532574
rect 171266 496658 171502 496894
rect 171586 496658 171822 496894
rect 171266 496338 171502 496574
rect 171586 496338 171822 496574
rect 192986 710362 193222 710598
rect 193306 710362 193542 710598
rect 192986 710042 193222 710278
rect 193306 710042 193542 710278
rect 189266 708442 189502 708678
rect 189586 708442 189822 708678
rect 189266 708122 189502 708358
rect 189586 708122 189822 708358
rect 185546 706522 185782 706758
rect 185866 706522 186102 706758
rect 185546 706202 185782 706438
rect 185866 706202 186102 706438
rect 174986 680378 175222 680614
rect 175306 680378 175542 680614
rect 174986 680058 175222 680294
rect 175306 680058 175542 680294
rect 174986 644378 175222 644614
rect 175306 644378 175542 644614
rect 174986 644058 175222 644294
rect 175306 644058 175542 644294
rect 174986 608378 175222 608614
rect 175306 608378 175542 608614
rect 174986 608058 175222 608294
rect 175306 608058 175542 608294
rect 174986 572378 175222 572614
rect 175306 572378 175542 572614
rect 174986 572058 175222 572294
rect 175306 572058 175542 572294
rect 174986 536378 175222 536614
rect 175306 536378 175542 536614
rect 174986 536058 175222 536294
rect 175306 536058 175542 536294
rect 174986 500378 175222 500614
rect 175306 500378 175542 500614
rect 174986 500058 175222 500294
rect 175306 500058 175542 500294
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 185546 690938 185782 691174
rect 185866 690938 186102 691174
rect 185546 690618 185782 690854
rect 185866 690618 186102 690854
rect 185546 654938 185782 655174
rect 185866 654938 186102 655174
rect 185546 654618 185782 654854
rect 185866 654618 186102 654854
rect 185546 618938 185782 619174
rect 185866 618938 186102 619174
rect 185546 618618 185782 618854
rect 185866 618618 186102 618854
rect 185546 582938 185782 583174
rect 185866 582938 186102 583174
rect 185546 582618 185782 582854
rect 185866 582618 186102 582854
rect 185546 546938 185782 547174
rect 185866 546938 186102 547174
rect 185546 546618 185782 546854
rect 185866 546618 186102 546854
rect 185546 510938 185782 511174
rect 185866 510938 186102 511174
rect 185546 510618 185782 510854
rect 185866 510618 186102 510854
rect 185546 474938 185782 475174
rect 185866 474938 186102 475174
rect 185546 474618 185782 474854
rect 185866 474618 186102 474854
rect 189266 694658 189502 694894
rect 189586 694658 189822 694894
rect 189266 694338 189502 694574
rect 189586 694338 189822 694574
rect 189266 658658 189502 658894
rect 189586 658658 189822 658894
rect 189266 658338 189502 658574
rect 189586 658338 189822 658574
rect 189266 622658 189502 622894
rect 189586 622658 189822 622894
rect 189266 622338 189502 622574
rect 189586 622338 189822 622574
rect 189266 586658 189502 586894
rect 189586 586658 189822 586894
rect 189266 586338 189502 586574
rect 189586 586338 189822 586574
rect 189266 550658 189502 550894
rect 189586 550658 189822 550894
rect 189266 550338 189502 550574
rect 189586 550338 189822 550574
rect 189266 514658 189502 514894
rect 189586 514658 189822 514894
rect 189266 514338 189502 514574
rect 189586 514338 189822 514574
rect 189266 478658 189502 478894
rect 189586 478658 189822 478894
rect 189266 478338 189502 478574
rect 189586 478338 189822 478574
rect 50328 453218 50564 453454
rect 50328 452898 50564 453134
rect 186056 453218 186292 453454
rect 186056 452898 186292 453134
rect 45266 442658 45502 442894
rect 45586 442658 45822 442894
rect 45266 442338 45502 442574
rect 45586 442338 45822 442574
rect 189266 442658 189502 442894
rect 189586 442658 189822 442894
rect 189266 442338 189502 442574
rect 189586 442338 189822 442574
rect 51008 435218 51244 435454
rect 51008 434898 51244 435134
rect 185376 435218 185612 435454
rect 185376 434898 185612 435134
rect 50328 417218 50564 417454
rect 50328 416898 50564 417134
rect 186056 417218 186292 417454
rect 186056 416898 186292 417134
rect 45266 406658 45502 406894
rect 45586 406658 45822 406894
rect 45266 406338 45502 406574
rect 45586 406338 45822 406574
rect 189266 406658 189502 406894
rect 189586 406658 189822 406894
rect 189266 406338 189502 406574
rect 189586 406338 189822 406574
rect 51008 399218 51244 399454
rect 51008 398898 51244 399134
rect 185376 399218 185612 399454
rect 185376 398898 185612 399134
rect 50328 381218 50564 381454
rect 50328 380898 50564 381134
rect 186056 381218 186292 381454
rect 186056 380898 186292 381134
rect 45266 370658 45502 370894
rect 45586 370658 45822 370894
rect 45266 370338 45502 370574
rect 45586 370338 45822 370574
rect 45266 334658 45502 334894
rect 45586 334658 45822 334894
rect 45266 334338 45502 334574
rect 45586 334338 45822 334574
rect 45266 298658 45502 298894
rect 45586 298658 45822 298894
rect 45266 298338 45502 298574
rect 45586 298338 45822 298574
rect 48986 374378 49222 374614
rect 49306 374378 49542 374614
rect 48986 374058 49222 374294
rect 49306 374058 49542 374294
rect 48986 338378 49222 338614
rect 49306 338378 49542 338614
rect 48986 338058 49222 338294
rect 49306 338058 49542 338294
rect 48986 302378 49222 302614
rect 49306 302378 49542 302614
rect 48986 302058 49222 302294
rect 49306 302058 49542 302294
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 59546 348938 59782 349174
rect 59866 348938 60102 349174
rect 59546 348618 59782 348854
rect 59866 348618 60102 348854
rect 59546 312938 59782 313174
rect 59866 312938 60102 313174
rect 59546 312618 59782 312854
rect 59866 312618 60102 312854
rect 63266 352658 63502 352894
rect 63586 352658 63822 352894
rect 63266 352338 63502 352574
rect 63586 352338 63822 352574
rect 63266 316658 63502 316894
rect 63586 316658 63822 316894
rect 63266 316338 63502 316574
rect 63586 316338 63822 316574
rect 66986 356378 67222 356614
rect 67306 356378 67542 356614
rect 66986 356058 67222 356294
rect 67306 356058 67542 356294
rect 66986 320378 67222 320614
rect 67306 320378 67542 320614
rect 66986 320058 67222 320294
rect 67306 320058 67542 320294
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 73826 327218 74062 327454
rect 74146 327218 74382 327454
rect 73826 326898 74062 327134
rect 74146 326898 74382 327134
rect 73826 291218 74062 291454
rect 74146 291218 74382 291454
rect 73826 290898 74062 291134
rect 74146 290898 74382 291134
rect 77546 366938 77782 367174
rect 77866 366938 78102 367174
rect 77546 366618 77782 366854
rect 77866 366618 78102 366854
rect 77546 330938 77782 331174
rect 77866 330938 78102 331174
rect 77546 330618 77782 330854
rect 77866 330618 78102 330854
rect 77546 294938 77782 295174
rect 77866 294938 78102 295174
rect 77546 294618 77782 294854
rect 77866 294618 78102 294854
rect 81266 370658 81502 370894
rect 81586 370658 81822 370894
rect 81266 370338 81502 370574
rect 81586 370338 81822 370574
rect 81266 334658 81502 334894
rect 81586 334658 81822 334894
rect 81266 334338 81502 334574
rect 81586 334338 81822 334574
rect 81266 298658 81502 298894
rect 81586 298658 81822 298894
rect 81266 298338 81502 298574
rect 81586 298338 81822 298574
rect 84986 374378 85222 374614
rect 85306 374378 85542 374614
rect 84986 374058 85222 374294
rect 85306 374058 85542 374294
rect 84986 338378 85222 338614
rect 85306 338378 85542 338614
rect 84986 338058 85222 338294
rect 85306 338058 85542 338294
rect 84986 302378 85222 302614
rect 85306 302378 85542 302614
rect 84986 302058 85222 302294
rect 85306 302058 85542 302294
rect 91826 345218 92062 345454
rect 92146 345218 92382 345454
rect 91826 344898 92062 345134
rect 92146 344898 92382 345134
rect 91826 309218 92062 309454
rect 92146 309218 92382 309454
rect 91826 308898 92062 309134
rect 92146 308898 92382 309134
rect 95546 348938 95782 349174
rect 95866 348938 96102 349174
rect 95546 348618 95782 348854
rect 95866 348618 96102 348854
rect 95546 312938 95782 313174
rect 95866 312938 96102 313174
rect 95546 312618 95782 312854
rect 95866 312618 96102 312854
rect 99266 352658 99502 352894
rect 99586 352658 99822 352894
rect 99266 352338 99502 352574
rect 99586 352338 99822 352574
rect 99266 316658 99502 316894
rect 99586 316658 99822 316894
rect 99266 316338 99502 316574
rect 99586 316338 99822 316574
rect 102986 356378 103222 356614
rect 103306 356378 103542 356614
rect 102986 356058 103222 356294
rect 103306 356058 103542 356294
rect 102986 320378 103222 320614
rect 103306 320378 103542 320614
rect 102986 320058 103222 320294
rect 103306 320058 103542 320294
rect 109826 363218 110062 363454
rect 110146 363218 110382 363454
rect 109826 362898 110062 363134
rect 110146 362898 110382 363134
rect 109826 327218 110062 327454
rect 110146 327218 110382 327454
rect 109826 326898 110062 327134
rect 110146 326898 110382 327134
rect 109826 291218 110062 291454
rect 110146 291218 110382 291454
rect 109826 290898 110062 291134
rect 110146 290898 110382 291134
rect 113546 366938 113782 367174
rect 113866 366938 114102 367174
rect 113546 366618 113782 366854
rect 113866 366618 114102 366854
rect 113546 330938 113782 331174
rect 113866 330938 114102 331174
rect 113546 330618 113782 330854
rect 113866 330618 114102 330854
rect 113546 294938 113782 295174
rect 113866 294938 114102 295174
rect 113546 294618 113782 294854
rect 113866 294618 114102 294854
rect 117266 370658 117502 370894
rect 117586 370658 117822 370894
rect 117266 370338 117502 370574
rect 117586 370338 117822 370574
rect 117266 334658 117502 334894
rect 117586 334658 117822 334894
rect 117266 334338 117502 334574
rect 117586 334338 117822 334574
rect 117266 298658 117502 298894
rect 117586 298658 117822 298894
rect 117266 298338 117502 298574
rect 117586 298338 117822 298574
rect 120986 374378 121222 374614
rect 121306 374378 121542 374614
rect 120986 374058 121222 374294
rect 121306 374058 121542 374294
rect 120986 338378 121222 338614
rect 121306 338378 121542 338614
rect 120986 338058 121222 338294
rect 121306 338058 121542 338294
rect 120986 302378 121222 302614
rect 121306 302378 121542 302614
rect 120986 302058 121222 302294
rect 121306 302058 121542 302294
rect 127826 345218 128062 345454
rect 128146 345218 128382 345454
rect 127826 344898 128062 345134
rect 128146 344898 128382 345134
rect 127826 309218 128062 309454
rect 128146 309218 128382 309454
rect 127826 308898 128062 309134
rect 128146 308898 128382 309134
rect 131546 348938 131782 349174
rect 131866 348938 132102 349174
rect 131546 348618 131782 348854
rect 131866 348618 132102 348854
rect 131546 312938 131782 313174
rect 131866 312938 132102 313174
rect 131546 312618 131782 312854
rect 131866 312618 132102 312854
rect 135266 352658 135502 352894
rect 135586 352658 135822 352894
rect 135266 352338 135502 352574
rect 135586 352338 135822 352574
rect 135266 316658 135502 316894
rect 135586 316658 135822 316894
rect 135266 316338 135502 316574
rect 135586 316338 135822 316574
rect 138986 356378 139222 356614
rect 139306 356378 139542 356614
rect 138986 356058 139222 356294
rect 139306 356058 139542 356294
rect 138986 320378 139222 320614
rect 139306 320378 139542 320614
rect 138986 320058 139222 320294
rect 139306 320058 139542 320294
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 145826 327218 146062 327454
rect 146146 327218 146382 327454
rect 145826 326898 146062 327134
rect 146146 326898 146382 327134
rect 145826 291218 146062 291454
rect 146146 291218 146382 291454
rect 145826 290898 146062 291134
rect 146146 290898 146382 291134
rect 149546 366938 149782 367174
rect 149866 366938 150102 367174
rect 149546 366618 149782 366854
rect 149866 366618 150102 366854
rect 149546 330938 149782 331174
rect 149866 330938 150102 331174
rect 149546 330618 149782 330854
rect 149866 330618 150102 330854
rect 149546 294938 149782 295174
rect 149866 294938 150102 295174
rect 149546 294618 149782 294854
rect 149866 294618 150102 294854
rect 153266 370658 153502 370894
rect 153586 370658 153822 370894
rect 153266 370338 153502 370574
rect 153586 370338 153822 370574
rect 153266 334658 153502 334894
rect 153586 334658 153822 334894
rect 153266 334338 153502 334574
rect 153586 334338 153822 334574
rect 153266 298658 153502 298894
rect 153586 298658 153822 298894
rect 153266 298338 153502 298574
rect 153586 298338 153822 298574
rect 156986 374378 157222 374614
rect 157306 374378 157542 374614
rect 156986 374058 157222 374294
rect 157306 374058 157542 374294
rect 156986 338378 157222 338614
rect 157306 338378 157542 338614
rect 156986 338058 157222 338294
rect 157306 338058 157542 338294
rect 156986 302378 157222 302614
rect 157306 302378 157542 302614
rect 156986 302058 157222 302294
rect 157306 302058 157542 302294
rect 163826 345218 164062 345454
rect 164146 345218 164382 345454
rect 163826 344898 164062 345134
rect 164146 344898 164382 345134
rect 163826 309218 164062 309454
rect 164146 309218 164382 309454
rect 163826 308898 164062 309134
rect 164146 308898 164382 309134
rect 167546 348938 167782 349174
rect 167866 348938 168102 349174
rect 167546 348618 167782 348854
rect 167866 348618 168102 348854
rect 167546 312938 167782 313174
rect 167866 312938 168102 313174
rect 167546 312618 167782 312854
rect 167866 312618 168102 312854
rect 171266 352658 171502 352894
rect 171586 352658 171822 352894
rect 171266 352338 171502 352574
rect 171586 352338 171822 352574
rect 171266 316658 171502 316894
rect 171586 316658 171822 316894
rect 171266 316338 171502 316574
rect 171586 316338 171822 316574
rect 174986 356378 175222 356614
rect 175306 356378 175542 356614
rect 174986 356058 175222 356294
rect 175306 356058 175542 356294
rect 174986 320378 175222 320614
rect 175306 320378 175542 320614
rect 174986 320058 175222 320294
rect 175306 320058 175542 320294
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 181826 327218 182062 327454
rect 182146 327218 182382 327454
rect 181826 326898 182062 327134
rect 182146 326898 182382 327134
rect 181826 291218 182062 291454
rect 182146 291218 182382 291454
rect 181826 290898 182062 291134
rect 182146 290898 182382 291134
rect 185546 366938 185782 367174
rect 185866 366938 186102 367174
rect 185546 366618 185782 366854
rect 185866 366618 186102 366854
rect 185546 330938 185782 331174
rect 185866 330938 186102 331174
rect 185546 330618 185782 330854
rect 185866 330618 186102 330854
rect 185546 294938 185782 295174
rect 185866 294938 186102 295174
rect 185546 294618 185782 294854
rect 185866 294618 186102 294854
rect 189266 370658 189502 370894
rect 189586 370658 189822 370894
rect 189266 370338 189502 370574
rect 189586 370338 189822 370574
rect 189266 334658 189502 334894
rect 189586 334658 189822 334894
rect 189266 334338 189502 334574
rect 189586 334338 189822 334574
rect 189266 298658 189502 298894
rect 189586 298658 189822 298894
rect 189266 298338 189502 298574
rect 189586 298338 189822 298574
rect 50328 273218 50564 273454
rect 50328 272898 50564 273134
rect 186056 273218 186292 273454
rect 186056 272898 186292 273134
rect 45266 262658 45502 262894
rect 45586 262658 45822 262894
rect 45266 262338 45502 262574
rect 45586 262338 45822 262574
rect 51008 255218 51244 255454
rect 51008 254898 51244 255134
rect 185376 255218 185612 255454
rect 185376 254898 185612 255134
rect 50328 237218 50564 237454
rect 50328 236898 50564 237134
rect 186056 237218 186292 237454
rect 186056 236898 186292 237134
rect 45266 226658 45502 226894
rect 45586 226658 45822 226894
rect 45266 226338 45502 226574
rect 45586 226338 45822 226574
rect 51008 219218 51244 219454
rect 51008 218898 51244 219134
rect 185376 219218 185612 219454
rect 185376 218898 185612 219134
rect 50328 201218 50564 201454
rect 50328 200898 50564 201134
rect 186056 201218 186292 201454
rect 186056 200898 186292 201134
rect 45266 190658 45502 190894
rect 45586 190658 45822 190894
rect 45266 190338 45502 190574
rect 45586 190338 45822 190574
rect 45266 154658 45502 154894
rect 45586 154658 45822 154894
rect 45266 154338 45502 154574
rect 45586 154338 45822 154574
rect 45266 118658 45502 118894
rect 45586 118658 45822 118894
rect 45266 118338 45502 118574
rect 45586 118338 45822 118574
rect 45266 82658 45502 82894
rect 45586 82658 45822 82894
rect 45266 82338 45502 82574
rect 45586 82338 45822 82574
rect 45266 46658 45502 46894
rect 45586 46658 45822 46894
rect 45266 46338 45502 46574
rect 45586 46338 45822 46574
rect 45266 10658 45502 10894
rect 45586 10658 45822 10894
rect 45266 10338 45502 10574
rect 45586 10338 45822 10574
rect 45266 -4422 45502 -4186
rect 45586 -4422 45822 -4186
rect 45266 -4742 45502 -4506
rect 45586 -4742 45822 -4506
rect 48986 194378 49222 194614
rect 49306 194378 49542 194614
rect 48986 194058 49222 194294
rect 49306 194058 49542 194294
rect 48986 158378 49222 158614
rect 49306 158378 49542 158614
rect 48986 158058 49222 158294
rect 49306 158058 49542 158294
rect 48986 122378 49222 122614
rect 49306 122378 49542 122614
rect 48986 122058 49222 122294
rect 49306 122058 49542 122294
rect 48986 86378 49222 86614
rect 49306 86378 49542 86614
rect 48986 86058 49222 86294
rect 49306 86058 49542 86294
rect 48986 50378 49222 50614
rect 49306 50378 49542 50614
rect 48986 50058 49222 50294
rect 49306 50058 49542 50294
rect 48986 14378 49222 14614
rect 49306 14378 49542 14614
rect 48986 14058 49222 14294
rect 49306 14058 49542 14294
rect 30986 -7302 31222 -7066
rect 31306 -7302 31542 -7066
rect 30986 -7622 31222 -7386
rect 31306 -7622 31542 -7386
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -1542 56062 -1306
rect 56146 -1542 56382 -1306
rect 55826 -1862 56062 -1626
rect 56146 -1862 56382 -1626
rect 59546 168938 59782 169174
rect 59866 168938 60102 169174
rect 59546 168618 59782 168854
rect 59866 168618 60102 168854
rect 59546 132938 59782 133174
rect 59866 132938 60102 133174
rect 59546 132618 59782 132854
rect 59866 132618 60102 132854
rect 59546 96938 59782 97174
rect 59866 96938 60102 97174
rect 59546 96618 59782 96854
rect 59866 96618 60102 96854
rect 59546 60938 59782 61174
rect 59866 60938 60102 61174
rect 59546 60618 59782 60854
rect 59866 60618 60102 60854
rect 59546 24938 59782 25174
rect 59866 24938 60102 25174
rect 59546 24618 59782 24854
rect 59866 24618 60102 24854
rect 59546 -3462 59782 -3226
rect 59866 -3462 60102 -3226
rect 59546 -3782 59782 -3546
rect 59866 -3782 60102 -3546
rect 63266 172658 63502 172894
rect 63586 172658 63822 172894
rect 63266 172338 63502 172574
rect 63586 172338 63822 172574
rect 63266 136658 63502 136894
rect 63586 136658 63822 136894
rect 63266 136338 63502 136574
rect 63586 136338 63822 136574
rect 63266 100658 63502 100894
rect 63586 100658 63822 100894
rect 63266 100338 63502 100574
rect 63586 100338 63822 100574
rect 63266 64658 63502 64894
rect 63586 64658 63822 64894
rect 63266 64338 63502 64574
rect 63586 64338 63822 64574
rect 63266 28658 63502 28894
rect 63586 28658 63822 28894
rect 63266 28338 63502 28574
rect 63586 28338 63822 28574
rect 63266 -5382 63502 -5146
rect 63586 -5382 63822 -5146
rect 63266 -5702 63502 -5466
rect 63586 -5702 63822 -5466
rect 66986 176378 67222 176614
rect 67306 176378 67542 176614
rect 66986 176058 67222 176294
rect 67306 176058 67542 176294
rect 66986 140378 67222 140614
rect 67306 140378 67542 140614
rect 66986 140058 67222 140294
rect 67306 140058 67542 140294
rect 66986 104378 67222 104614
rect 67306 104378 67542 104614
rect 66986 104058 67222 104294
rect 67306 104058 67542 104294
rect 66986 68378 67222 68614
rect 67306 68378 67542 68614
rect 66986 68058 67222 68294
rect 67306 68058 67542 68294
rect 66986 32378 67222 32614
rect 67306 32378 67542 32614
rect 66986 32058 67222 32294
rect 67306 32058 67542 32294
rect 48986 -6342 49222 -6106
rect 49306 -6342 49542 -6106
rect 48986 -6662 49222 -6426
rect 49306 -6662 49542 -6426
rect 73826 183218 74062 183454
rect 74146 183218 74382 183454
rect 73826 182898 74062 183134
rect 74146 182898 74382 183134
rect 73826 147218 74062 147454
rect 74146 147218 74382 147454
rect 73826 146898 74062 147134
rect 74146 146898 74382 147134
rect 73826 111218 74062 111454
rect 74146 111218 74382 111454
rect 73826 110898 74062 111134
rect 74146 110898 74382 111134
rect 73826 75218 74062 75454
rect 74146 75218 74382 75454
rect 73826 74898 74062 75134
rect 74146 74898 74382 75134
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 186938 77782 187174
rect 77866 186938 78102 187174
rect 77546 186618 77782 186854
rect 77866 186618 78102 186854
rect 77546 150938 77782 151174
rect 77866 150938 78102 151174
rect 77546 150618 77782 150854
rect 77866 150618 78102 150854
rect 77546 114938 77782 115174
rect 77866 114938 78102 115174
rect 77546 114618 77782 114854
rect 77866 114618 78102 114854
rect 77546 78938 77782 79174
rect 77866 78938 78102 79174
rect 77546 78618 77782 78854
rect 77866 78618 78102 78854
rect 77546 42938 77782 43174
rect 77866 42938 78102 43174
rect 77546 42618 77782 42854
rect 77866 42618 78102 42854
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -2502 77782 -2266
rect 77866 -2502 78102 -2266
rect 77546 -2822 77782 -2586
rect 77866 -2822 78102 -2586
rect 81266 190658 81502 190894
rect 81586 190658 81822 190894
rect 81266 190338 81502 190574
rect 81586 190338 81822 190574
rect 81266 154658 81502 154894
rect 81586 154658 81822 154894
rect 81266 154338 81502 154574
rect 81586 154338 81822 154574
rect 81266 118658 81502 118894
rect 81586 118658 81822 118894
rect 81266 118338 81502 118574
rect 81586 118338 81822 118574
rect 81266 82658 81502 82894
rect 81586 82658 81822 82894
rect 81266 82338 81502 82574
rect 81586 82338 81822 82574
rect 81266 46658 81502 46894
rect 81586 46658 81822 46894
rect 81266 46338 81502 46574
rect 81586 46338 81822 46574
rect 81266 10658 81502 10894
rect 81586 10658 81822 10894
rect 81266 10338 81502 10574
rect 81586 10338 81822 10574
rect 81266 -4422 81502 -4186
rect 81586 -4422 81822 -4186
rect 81266 -4742 81502 -4506
rect 81586 -4742 81822 -4506
rect 84986 194378 85222 194614
rect 85306 194378 85542 194614
rect 84986 194058 85222 194294
rect 85306 194058 85542 194294
rect 84986 158378 85222 158614
rect 85306 158378 85542 158614
rect 84986 158058 85222 158294
rect 85306 158058 85542 158294
rect 84986 122378 85222 122614
rect 85306 122378 85542 122614
rect 84986 122058 85222 122294
rect 85306 122058 85542 122294
rect 84986 86378 85222 86614
rect 85306 86378 85542 86614
rect 84986 86058 85222 86294
rect 85306 86058 85542 86294
rect 84986 50378 85222 50614
rect 85306 50378 85542 50614
rect 84986 50058 85222 50294
rect 85306 50058 85542 50294
rect 84986 14378 85222 14614
rect 85306 14378 85542 14614
rect 84986 14058 85222 14294
rect 85306 14058 85542 14294
rect 66986 -7302 67222 -7066
rect 67306 -7302 67542 -7066
rect 66986 -7622 67222 -7386
rect 67306 -7622 67542 -7386
rect 91826 165218 92062 165454
rect 92146 165218 92382 165454
rect 91826 164898 92062 165134
rect 92146 164898 92382 165134
rect 91826 129218 92062 129454
rect 92146 129218 92382 129454
rect 91826 128898 92062 129134
rect 92146 128898 92382 129134
rect 91826 93218 92062 93454
rect 92146 93218 92382 93454
rect 91826 92898 92062 93134
rect 92146 92898 92382 93134
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -1542 92062 -1306
rect 92146 -1542 92382 -1306
rect 91826 -1862 92062 -1626
rect 92146 -1862 92382 -1626
rect 95546 168938 95782 169174
rect 95866 168938 96102 169174
rect 95546 168618 95782 168854
rect 95866 168618 96102 168854
rect 95546 132938 95782 133174
rect 95866 132938 96102 133174
rect 95546 132618 95782 132854
rect 95866 132618 96102 132854
rect 95546 96938 95782 97174
rect 95866 96938 96102 97174
rect 95546 96618 95782 96854
rect 95866 96618 96102 96854
rect 95546 60938 95782 61174
rect 95866 60938 96102 61174
rect 95546 60618 95782 60854
rect 95866 60618 96102 60854
rect 95546 24938 95782 25174
rect 95866 24938 96102 25174
rect 95546 24618 95782 24854
rect 95866 24618 96102 24854
rect 95546 -3462 95782 -3226
rect 95866 -3462 96102 -3226
rect 95546 -3782 95782 -3546
rect 95866 -3782 96102 -3546
rect 99266 172658 99502 172894
rect 99586 172658 99822 172894
rect 99266 172338 99502 172574
rect 99586 172338 99822 172574
rect 99266 136658 99502 136894
rect 99586 136658 99822 136894
rect 99266 136338 99502 136574
rect 99586 136338 99822 136574
rect 99266 100658 99502 100894
rect 99586 100658 99822 100894
rect 99266 100338 99502 100574
rect 99586 100338 99822 100574
rect 99266 64658 99502 64894
rect 99586 64658 99822 64894
rect 99266 64338 99502 64574
rect 99586 64338 99822 64574
rect 99266 28658 99502 28894
rect 99586 28658 99822 28894
rect 99266 28338 99502 28574
rect 99586 28338 99822 28574
rect 99266 -5382 99502 -5146
rect 99586 -5382 99822 -5146
rect 99266 -5702 99502 -5466
rect 99586 -5702 99822 -5466
rect 102986 176378 103222 176614
rect 103306 176378 103542 176614
rect 102986 176058 103222 176294
rect 103306 176058 103542 176294
rect 102986 140378 103222 140614
rect 103306 140378 103542 140614
rect 102986 140058 103222 140294
rect 103306 140058 103542 140294
rect 102986 104378 103222 104614
rect 103306 104378 103542 104614
rect 102986 104058 103222 104294
rect 103306 104058 103542 104294
rect 102986 68378 103222 68614
rect 103306 68378 103542 68614
rect 102986 68058 103222 68294
rect 103306 68058 103542 68294
rect 102986 32378 103222 32614
rect 103306 32378 103542 32614
rect 102986 32058 103222 32294
rect 103306 32058 103542 32294
rect 84986 -6342 85222 -6106
rect 85306 -6342 85542 -6106
rect 84986 -6662 85222 -6426
rect 85306 -6662 85542 -6426
rect 109826 183218 110062 183454
rect 110146 183218 110382 183454
rect 109826 182898 110062 183134
rect 110146 182898 110382 183134
rect 109826 147218 110062 147454
rect 110146 147218 110382 147454
rect 109826 146898 110062 147134
rect 110146 146898 110382 147134
rect 109826 111218 110062 111454
rect 110146 111218 110382 111454
rect 109826 110898 110062 111134
rect 110146 110898 110382 111134
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 186938 113782 187174
rect 113866 186938 114102 187174
rect 113546 186618 113782 186854
rect 113866 186618 114102 186854
rect 113546 150938 113782 151174
rect 113866 150938 114102 151174
rect 113546 150618 113782 150854
rect 113866 150618 114102 150854
rect 113546 114938 113782 115174
rect 113866 114938 114102 115174
rect 113546 114618 113782 114854
rect 113866 114618 114102 114854
rect 113546 78938 113782 79174
rect 113866 78938 114102 79174
rect 113546 78618 113782 78854
rect 113866 78618 114102 78854
rect 113546 42938 113782 43174
rect 113866 42938 114102 43174
rect 113546 42618 113782 42854
rect 113866 42618 114102 42854
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 113546 -2502 113782 -2266
rect 113866 -2502 114102 -2266
rect 113546 -2822 113782 -2586
rect 113866 -2822 114102 -2586
rect 117266 190658 117502 190894
rect 117586 190658 117822 190894
rect 117266 190338 117502 190574
rect 117586 190338 117822 190574
rect 117266 154658 117502 154894
rect 117586 154658 117822 154894
rect 117266 154338 117502 154574
rect 117586 154338 117822 154574
rect 117266 118658 117502 118894
rect 117586 118658 117822 118894
rect 117266 118338 117502 118574
rect 117586 118338 117822 118574
rect 117266 82658 117502 82894
rect 117586 82658 117822 82894
rect 117266 82338 117502 82574
rect 117586 82338 117822 82574
rect 117266 46658 117502 46894
rect 117586 46658 117822 46894
rect 117266 46338 117502 46574
rect 117586 46338 117822 46574
rect 117266 10658 117502 10894
rect 117586 10658 117822 10894
rect 117266 10338 117502 10574
rect 117586 10338 117822 10574
rect 117266 -4422 117502 -4186
rect 117586 -4422 117822 -4186
rect 117266 -4742 117502 -4506
rect 117586 -4742 117822 -4506
rect 120986 194378 121222 194614
rect 121306 194378 121542 194614
rect 120986 194058 121222 194294
rect 121306 194058 121542 194294
rect 120986 158378 121222 158614
rect 121306 158378 121542 158614
rect 120986 158058 121222 158294
rect 121306 158058 121542 158294
rect 120986 122378 121222 122614
rect 121306 122378 121542 122614
rect 120986 122058 121222 122294
rect 121306 122058 121542 122294
rect 120986 86378 121222 86614
rect 121306 86378 121542 86614
rect 120986 86058 121222 86294
rect 121306 86058 121542 86294
rect 120986 50378 121222 50614
rect 121306 50378 121542 50614
rect 120986 50058 121222 50294
rect 121306 50058 121542 50294
rect 120986 14378 121222 14614
rect 121306 14378 121542 14614
rect 120986 14058 121222 14294
rect 121306 14058 121542 14294
rect 102986 -7302 103222 -7066
rect 103306 -7302 103542 -7066
rect 102986 -7622 103222 -7386
rect 103306 -7622 103542 -7386
rect 127826 165218 128062 165454
rect 128146 165218 128382 165454
rect 127826 164898 128062 165134
rect 128146 164898 128382 165134
rect 127826 129218 128062 129454
rect 128146 129218 128382 129454
rect 127826 128898 128062 129134
rect 128146 128898 128382 129134
rect 127826 93218 128062 93454
rect 128146 93218 128382 93454
rect 127826 92898 128062 93134
rect 128146 92898 128382 93134
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -1542 128062 -1306
rect 128146 -1542 128382 -1306
rect 127826 -1862 128062 -1626
rect 128146 -1862 128382 -1626
rect 131546 168938 131782 169174
rect 131866 168938 132102 169174
rect 131546 168618 131782 168854
rect 131866 168618 132102 168854
rect 131546 132938 131782 133174
rect 131866 132938 132102 133174
rect 131546 132618 131782 132854
rect 131866 132618 132102 132854
rect 131546 96938 131782 97174
rect 131866 96938 132102 97174
rect 131546 96618 131782 96854
rect 131866 96618 132102 96854
rect 131546 60938 131782 61174
rect 131866 60938 132102 61174
rect 131546 60618 131782 60854
rect 131866 60618 132102 60854
rect 131546 24938 131782 25174
rect 131866 24938 132102 25174
rect 131546 24618 131782 24854
rect 131866 24618 132102 24854
rect 131546 -3462 131782 -3226
rect 131866 -3462 132102 -3226
rect 131546 -3782 131782 -3546
rect 131866 -3782 132102 -3546
rect 135266 172658 135502 172894
rect 135586 172658 135822 172894
rect 135266 172338 135502 172574
rect 135586 172338 135822 172574
rect 135266 136658 135502 136894
rect 135586 136658 135822 136894
rect 135266 136338 135502 136574
rect 135586 136338 135822 136574
rect 135266 100658 135502 100894
rect 135586 100658 135822 100894
rect 135266 100338 135502 100574
rect 135586 100338 135822 100574
rect 135266 64658 135502 64894
rect 135586 64658 135822 64894
rect 135266 64338 135502 64574
rect 135586 64338 135822 64574
rect 135266 28658 135502 28894
rect 135586 28658 135822 28894
rect 135266 28338 135502 28574
rect 135586 28338 135822 28574
rect 135266 -5382 135502 -5146
rect 135586 -5382 135822 -5146
rect 135266 -5702 135502 -5466
rect 135586 -5702 135822 -5466
rect 138986 176378 139222 176614
rect 139306 176378 139542 176614
rect 138986 176058 139222 176294
rect 139306 176058 139542 176294
rect 138986 140378 139222 140614
rect 139306 140378 139542 140614
rect 138986 140058 139222 140294
rect 139306 140058 139542 140294
rect 138986 104378 139222 104614
rect 139306 104378 139542 104614
rect 138986 104058 139222 104294
rect 139306 104058 139542 104294
rect 138986 68378 139222 68614
rect 139306 68378 139542 68614
rect 138986 68058 139222 68294
rect 139306 68058 139542 68294
rect 138986 32378 139222 32614
rect 139306 32378 139542 32614
rect 138986 32058 139222 32294
rect 139306 32058 139542 32294
rect 120986 -6342 121222 -6106
rect 121306 -6342 121542 -6106
rect 120986 -6662 121222 -6426
rect 121306 -6662 121542 -6426
rect 145826 183218 146062 183454
rect 146146 183218 146382 183454
rect 145826 182898 146062 183134
rect 146146 182898 146382 183134
rect 145826 147218 146062 147454
rect 146146 147218 146382 147454
rect 145826 146898 146062 147134
rect 146146 146898 146382 147134
rect 145826 111218 146062 111454
rect 146146 111218 146382 111454
rect 145826 110898 146062 111134
rect 146146 110898 146382 111134
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 186938 149782 187174
rect 149866 186938 150102 187174
rect 149546 186618 149782 186854
rect 149866 186618 150102 186854
rect 149546 150938 149782 151174
rect 149866 150938 150102 151174
rect 149546 150618 149782 150854
rect 149866 150618 150102 150854
rect 149546 114938 149782 115174
rect 149866 114938 150102 115174
rect 149546 114618 149782 114854
rect 149866 114618 150102 114854
rect 149546 78938 149782 79174
rect 149866 78938 150102 79174
rect 149546 78618 149782 78854
rect 149866 78618 150102 78854
rect 149546 42938 149782 43174
rect 149866 42938 150102 43174
rect 149546 42618 149782 42854
rect 149866 42618 150102 42854
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 149546 -2502 149782 -2266
rect 149866 -2502 150102 -2266
rect 149546 -2822 149782 -2586
rect 149866 -2822 150102 -2586
rect 153266 190658 153502 190894
rect 153586 190658 153822 190894
rect 153266 190338 153502 190574
rect 153586 190338 153822 190574
rect 153266 154658 153502 154894
rect 153586 154658 153822 154894
rect 153266 154338 153502 154574
rect 153586 154338 153822 154574
rect 153266 118658 153502 118894
rect 153586 118658 153822 118894
rect 153266 118338 153502 118574
rect 153586 118338 153822 118574
rect 153266 82658 153502 82894
rect 153586 82658 153822 82894
rect 153266 82338 153502 82574
rect 153586 82338 153822 82574
rect 153266 46658 153502 46894
rect 153586 46658 153822 46894
rect 153266 46338 153502 46574
rect 153586 46338 153822 46574
rect 153266 10658 153502 10894
rect 153586 10658 153822 10894
rect 153266 10338 153502 10574
rect 153586 10338 153822 10574
rect 153266 -4422 153502 -4186
rect 153586 -4422 153822 -4186
rect 153266 -4742 153502 -4506
rect 153586 -4742 153822 -4506
rect 156986 194378 157222 194614
rect 157306 194378 157542 194614
rect 156986 194058 157222 194294
rect 157306 194058 157542 194294
rect 156986 158378 157222 158614
rect 157306 158378 157542 158614
rect 156986 158058 157222 158294
rect 157306 158058 157542 158294
rect 156986 122378 157222 122614
rect 157306 122378 157542 122614
rect 156986 122058 157222 122294
rect 157306 122058 157542 122294
rect 156986 86378 157222 86614
rect 157306 86378 157542 86614
rect 156986 86058 157222 86294
rect 157306 86058 157542 86294
rect 156986 50378 157222 50614
rect 157306 50378 157542 50614
rect 156986 50058 157222 50294
rect 157306 50058 157542 50294
rect 156986 14378 157222 14614
rect 157306 14378 157542 14614
rect 156986 14058 157222 14294
rect 157306 14058 157542 14294
rect 138986 -7302 139222 -7066
rect 139306 -7302 139542 -7066
rect 138986 -7622 139222 -7386
rect 139306 -7622 139542 -7386
rect 163826 165218 164062 165454
rect 164146 165218 164382 165454
rect 163826 164898 164062 165134
rect 164146 164898 164382 165134
rect 163826 129218 164062 129454
rect 164146 129218 164382 129454
rect 163826 128898 164062 129134
rect 164146 128898 164382 129134
rect 163826 93218 164062 93454
rect 164146 93218 164382 93454
rect 163826 92898 164062 93134
rect 164146 92898 164382 93134
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -1542 164062 -1306
rect 164146 -1542 164382 -1306
rect 163826 -1862 164062 -1626
rect 164146 -1862 164382 -1626
rect 167546 168938 167782 169174
rect 167866 168938 168102 169174
rect 167546 168618 167782 168854
rect 167866 168618 168102 168854
rect 167546 132938 167782 133174
rect 167866 132938 168102 133174
rect 167546 132618 167782 132854
rect 167866 132618 168102 132854
rect 167546 96938 167782 97174
rect 167866 96938 168102 97174
rect 167546 96618 167782 96854
rect 167866 96618 168102 96854
rect 167546 60938 167782 61174
rect 167866 60938 168102 61174
rect 167546 60618 167782 60854
rect 167866 60618 168102 60854
rect 167546 24938 167782 25174
rect 167866 24938 168102 25174
rect 167546 24618 167782 24854
rect 167866 24618 168102 24854
rect 167546 -3462 167782 -3226
rect 167866 -3462 168102 -3226
rect 167546 -3782 167782 -3546
rect 167866 -3782 168102 -3546
rect 171266 172658 171502 172894
rect 171586 172658 171822 172894
rect 171266 172338 171502 172574
rect 171586 172338 171822 172574
rect 171266 136658 171502 136894
rect 171586 136658 171822 136894
rect 171266 136338 171502 136574
rect 171586 136338 171822 136574
rect 171266 100658 171502 100894
rect 171586 100658 171822 100894
rect 171266 100338 171502 100574
rect 171586 100338 171822 100574
rect 171266 64658 171502 64894
rect 171586 64658 171822 64894
rect 171266 64338 171502 64574
rect 171586 64338 171822 64574
rect 171266 28658 171502 28894
rect 171586 28658 171822 28894
rect 171266 28338 171502 28574
rect 171586 28338 171822 28574
rect 171266 -5382 171502 -5146
rect 171586 -5382 171822 -5146
rect 171266 -5702 171502 -5466
rect 171586 -5702 171822 -5466
rect 174986 176378 175222 176614
rect 175306 176378 175542 176614
rect 174986 176058 175222 176294
rect 175306 176058 175542 176294
rect 174986 140378 175222 140614
rect 175306 140378 175542 140614
rect 174986 140058 175222 140294
rect 175306 140058 175542 140294
rect 174986 104378 175222 104614
rect 175306 104378 175542 104614
rect 174986 104058 175222 104294
rect 175306 104058 175542 104294
rect 174986 68378 175222 68614
rect 175306 68378 175542 68614
rect 174986 68058 175222 68294
rect 175306 68058 175542 68294
rect 174986 32378 175222 32614
rect 175306 32378 175542 32614
rect 174986 32058 175222 32294
rect 175306 32058 175542 32294
rect 156986 -6342 157222 -6106
rect 157306 -6342 157542 -6106
rect 156986 -6662 157222 -6426
rect 157306 -6662 157542 -6426
rect 181826 183218 182062 183454
rect 182146 183218 182382 183454
rect 181826 182898 182062 183134
rect 182146 182898 182382 183134
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 181826 111218 182062 111454
rect 182146 111218 182382 111454
rect 181826 110898 182062 111134
rect 182146 110898 182382 111134
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 189266 262658 189502 262894
rect 189586 262658 189822 262894
rect 189266 262338 189502 262574
rect 189586 262338 189822 262574
rect 189266 226658 189502 226894
rect 189586 226658 189822 226894
rect 189266 226338 189502 226574
rect 189586 226338 189822 226574
rect 185546 186938 185782 187174
rect 185866 186938 186102 187174
rect 185546 186618 185782 186854
rect 185866 186618 186102 186854
rect 185546 150938 185782 151174
rect 185866 150938 186102 151174
rect 185546 150618 185782 150854
rect 185866 150618 186102 150854
rect 185546 114938 185782 115174
rect 185866 114938 186102 115174
rect 185546 114618 185782 114854
rect 185866 114618 186102 114854
rect 185546 78938 185782 79174
rect 185866 78938 186102 79174
rect 185546 78618 185782 78854
rect 185866 78618 186102 78854
rect 185546 42938 185782 43174
rect 185866 42938 186102 43174
rect 185546 42618 185782 42854
rect 185866 42618 186102 42854
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 185546 -2502 185782 -2266
rect 185866 -2502 186102 -2266
rect 185546 -2822 185782 -2586
rect 185866 -2822 186102 -2586
rect 189266 190658 189502 190894
rect 189586 190658 189822 190894
rect 189266 190338 189502 190574
rect 189586 190338 189822 190574
rect 189266 154658 189502 154894
rect 189586 154658 189822 154894
rect 189266 154338 189502 154574
rect 189586 154338 189822 154574
rect 189266 118658 189502 118894
rect 189586 118658 189822 118894
rect 189266 118338 189502 118574
rect 189586 118338 189822 118574
rect 189266 82658 189502 82894
rect 189586 82658 189822 82894
rect 189266 82338 189502 82574
rect 189586 82338 189822 82574
rect 189266 46658 189502 46894
rect 189586 46658 189822 46894
rect 189266 46338 189502 46574
rect 189586 46338 189822 46574
rect 189266 10658 189502 10894
rect 189586 10658 189822 10894
rect 189266 10338 189502 10574
rect 189586 10338 189822 10574
rect 189266 -4422 189502 -4186
rect 189586 -4422 189822 -4186
rect 189266 -4742 189502 -4506
rect 189586 -4742 189822 -4506
rect 210986 711322 211222 711558
rect 211306 711322 211542 711558
rect 210986 711002 211222 711238
rect 211306 711002 211542 711238
rect 207266 709402 207502 709638
rect 207586 709402 207822 709638
rect 207266 709082 207502 709318
rect 207586 709082 207822 709318
rect 203546 707482 203782 707718
rect 203866 707482 204102 707718
rect 203546 707162 203782 707398
rect 203866 707162 204102 707398
rect 192986 698378 193222 698614
rect 193306 698378 193542 698614
rect 192986 698058 193222 698294
rect 193306 698058 193542 698294
rect 192986 662378 193222 662614
rect 193306 662378 193542 662614
rect 192986 662058 193222 662294
rect 193306 662058 193542 662294
rect 192986 626378 193222 626614
rect 193306 626378 193542 626614
rect 192986 626058 193222 626294
rect 193306 626058 193542 626294
rect 192986 590378 193222 590614
rect 193306 590378 193542 590614
rect 192986 590058 193222 590294
rect 193306 590058 193542 590294
rect 192986 554378 193222 554614
rect 193306 554378 193542 554614
rect 192986 554058 193222 554294
rect 193306 554058 193542 554294
rect 192986 518378 193222 518614
rect 193306 518378 193542 518614
rect 192986 518058 193222 518294
rect 193306 518058 193542 518294
rect 192986 482378 193222 482614
rect 193306 482378 193542 482614
rect 192986 482058 193222 482294
rect 193306 482058 193542 482294
rect 192986 446378 193222 446614
rect 193306 446378 193542 446614
rect 192986 446058 193222 446294
rect 193306 446058 193542 446294
rect 192986 410378 193222 410614
rect 193306 410378 193542 410614
rect 192986 410058 193222 410294
rect 193306 410058 193542 410294
rect 192986 374378 193222 374614
rect 193306 374378 193542 374614
rect 192986 374058 193222 374294
rect 193306 374058 193542 374294
rect 192986 338378 193222 338614
rect 193306 338378 193542 338614
rect 192986 338058 193222 338294
rect 193306 338058 193542 338294
rect 192986 302378 193222 302614
rect 193306 302378 193542 302614
rect 192986 302058 193222 302294
rect 193306 302058 193542 302294
rect 192986 266378 193222 266614
rect 193306 266378 193542 266614
rect 192986 266058 193222 266294
rect 193306 266058 193542 266294
rect 192986 230378 193222 230614
rect 193306 230378 193542 230614
rect 192986 230058 193222 230294
rect 193306 230058 193542 230294
rect 192986 194378 193222 194614
rect 193306 194378 193542 194614
rect 192986 194058 193222 194294
rect 193306 194058 193542 194294
rect 192986 158378 193222 158614
rect 193306 158378 193542 158614
rect 192986 158058 193222 158294
rect 193306 158058 193542 158294
rect 192986 122378 193222 122614
rect 193306 122378 193542 122614
rect 192986 122058 193222 122294
rect 193306 122058 193542 122294
rect 192986 86378 193222 86614
rect 193306 86378 193542 86614
rect 192986 86058 193222 86294
rect 193306 86058 193542 86294
rect 192986 50378 193222 50614
rect 193306 50378 193542 50614
rect 192986 50058 193222 50294
rect 193306 50058 193542 50294
rect 192986 14378 193222 14614
rect 193306 14378 193542 14614
rect 192986 14058 193222 14294
rect 193306 14058 193542 14294
rect 174986 -7302 175222 -7066
rect 175306 -7302 175542 -7066
rect 174986 -7622 175222 -7386
rect 175306 -7622 175542 -7386
rect 199826 705562 200062 705798
rect 200146 705562 200382 705798
rect 199826 705242 200062 705478
rect 200146 705242 200382 705478
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 199826 561218 200062 561454
rect 200146 561218 200382 561454
rect 199826 560898 200062 561134
rect 200146 560898 200382 561134
rect 199826 525218 200062 525454
rect 200146 525218 200382 525454
rect 199826 524898 200062 525134
rect 200146 524898 200382 525134
rect 199826 489218 200062 489454
rect 200146 489218 200382 489454
rect 199826 488898 200062 489134
rect 200146 488898 200382 489134
rect 199826 453218 200062 453454
rect 200146 453218 200382 453454
rect 199826 452898 200062 453134
rect 200146 452898 200382 453134
rect 199826 417218 200062 417454
rect 200146 417218 200382 417454
rect 199826 416898 200062 417134
rect 200146 416898 200382 417134
rect 199826 381218 200062 381454
rect 200146 381218 200382 381454
rect 199826 380898 200062 381134
rect 200146 380898 200382 381134
rect 199826 345218 200062 345454
rect 200146 345218 200382 345454
rect 199826 344898 200062 345134
rect 200146 344898 200382 345134
rect 199826 309218 200062 309454
rect 200146 309218 200382 309454
rect 199826 308898 200062 309134
rect 200146 308898 200382 309134
rect 199826 273218 200062 273454
rect 200146 273218 200382 273454
rect 199826 272898 200062 273134
rect 200146 272898 200382 273134
rect 199826 237218 200062 237454
rect 200146 237218 200382 237454
rect 199826 236898 200062 237134
rect 200146 236898 200382 237134
rect 199826 201218 200062 201454
rect 200146 201218 200382 201454
rect 199826 200898 200062 201134
rect 200146 200898 200382 201134
rect 199826 165218 200062 165454
rect 200146 165218 200382 165454
rect 199826 164898 200062 165134
rect 200146 164898 200382 165134
rect 199826 129218 200062 129454
rect 200146 129218 200382 129454
rect 199826 128898 200062 129134
rect 200146 128898 200382 129134
rect 199826 93218 200062 93454
rect 200146 93218 200382 93454
rect 199826 92898 200062 93134
rect 200146 92898 200382 93134
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -1542 200062 -1306
rect 200146 -1542 200382 -1306
rect 199826 -1862 200062 -1626
rect 200146 -1862 200382 -1626
rect 203546 672938 203782 673174
rect 203866 672938 204102 673174
rect 203546 672618 203782 672854
rect 203866 672618 204102 672854
rect 203546 636938 203782 637174
rect 203866 636938 204102 637174
rect 203546 636618 203782 636854
rect 203866 636618 204102 636854
rect 203546 600938 203782 601174
rect 203866 600938 204102 601174
rect 203546 600618 203782 600854
rect 203866 600618 204102 600854
rect 203546 564938 203782 565174
rect 203866 564938 204102 565174
rect 203546 564618 203782 564854
rect 203866 564618 204102 564854
rect 203546 528938 203782 529174
rect 203866 528938 204102 529174
rect 203546 528618 203782 528854
rect 203866 528618 204102 528854
rect 203546 492938 203782 493174
rect 203866 492938 204102 493174
rect 203546 492618 203782 492854
rect 203866 492618 204102 492854
rect 203546 456938 203782 457174
rect 203866 456938 204102 457174
rect 203546 456618 203782 456854
rect 203866 456618 204102 456854
rect 203546 420938 203782 421174
rect 203866 420938 204102 421174
rect 203546 420618 203782 420854
rect 203866 420618 204102 420854
rect 203546 384938 203782 385174
rect 203866 384938 204102 385174
rect 203546 384618 203782 384854
rect 203866 384618 204102 384854
rect 203546 348938 203782 349174
rect 203866 348938 204102 349174
rect 203546 348618 203782 348854
rect 203866 348618 204102 348854
rect 203546 312938 203782 313174
rect 203866 312938 204102 313174
rect 203546 312618 203782 312854
rect 203866 312618 204102 312854
rect 203546 276938 203782 277174
rect 203866 276938 204102 277174
rect 203546 276618 203782 276854
rect 203866 276618 204102 276854
rect 203546 240938 203782 241174
rect 203866 240938 204102 241174
rect 203546 240618 203782 240854
rect 203866 240618 204102 240854
rect 203546 204938 203782 205174
rect 203866 204938 204102 205174
rect 203546 204618 203782 204854
rect 203866 204618 204102 204854
rect 203546 168938 203782 169174
rect 203866 168938 204102 169174
rect 203546 168618 203782 168854
rect 203866 168618 204102 168854
rect 203546 132938 203782 133174
rect 203866 132938 204102 133174
rect 203546 132618 203782 132854
rect 203866 132618 204102 132854
rect 203546 96938 203782 97174
rect 203866 96938 204102 97174
rect 203546 96618 203782 96854
rect 203866 96618 204102 96854
rect 203546 60938 203782 61174
rect 203866 60938 204102 61174
rect 203546 60618 203782 60854
rect 203866 60618 204102 60854
rect 203546 24938 203782 25174
rect 203866 24938 204102 25174
rect 203546 24618 203782 24854
rect 203866 24618 204102 24854
rect 203546 -3462 203782 -3226
rect 203866 -3462 204102 -3226
rect 203546 -3782 203782 -3546
rect 203866 -3782 204102 -3546
rect 207266 676658 207502 676894
rect 207586 676658 207822 676894
rect 207266 676338 207502 676574
rect 207586 676338 207822 676574
rect 207266 640658 207502 640894
rect 207586 640658 207822 640894
rect 207266 640338 207502 640574
rect 207586 640338 207822 640574
rect 207266 604658 207502 604894
rect 207586 604658 207822 604894
rect 207266 604338 207502 604574
rect 207586 604338 207822 604574
rect 207266 568658 207502 568894
rect 207586 568658 207822 568894
rect 207266 568338 207502 568574
rect 207586 568338 207822 568574
rect 207266 532658 207502 532894
rect 207586 532658 207822 532894
rect 207266 532338 207502 532574
rect 207586 532338 207822 532574
rect 207266 496658 207502 496894
rect 207586 496658 207822 496894
rect 207266 496338 207502 496574
rect 207586 496338 207822 496574
rect 207266 460658 207502 460894
rect 207586 460658 207822 460894
rect 207266 460338 207502 460574
rect 207586 460338 207822 460574
rect 207266 424658 207502 424894
rect 207586 424658 207822 424894
rect 207266 424338 207502 424574
rect 207586 424338 207822 424574
rect 207266 388658 207502 388894
rect 207586 388658 207822 388894
rect 207266 388338 207502 388574
rect 207586 388338 207822 388574
rect 207266 352658 207502 352894
rect 207586 352658 207822 352894
rect 207266 352338 207502 352574
rect 207586 352338 207822 352574
rect 207266 316658 207502 316894
rect 207586 316658 207822 316894
rect 207266 316338 207502 316574
rect 207586 316338 207822 316574
rect 207266 280658 207502 280894
rect 207586 280658 207822 280894
rect 207266 280338 207502 280574
rect 207586 280338 207822 280574
rect 207266 244658 207502 244894
rect 207586 244658 207822 244894
rect 207266 244338 207502 244574
rect 207586 244338 207822 244574
rect 207266 208658 207502 208894
rect 207586 208658 207822 208894
rect 207266 208338 207502 208574
rect 207586 208338 207822 208574
rect 207266 172658 207502 172894
rect 207586 172658 207822 172894
rect 207266 172338 207502 172574
rect 207586 172338 207822 172574
rect 207266 136658 207502 136894
rect 207586 136658 207822 136894
rect 207266 136338 207502 136574
rect 207586 136338 207822 136574
rect 207266 100658 207502 100894
rect 207586 100658 207822 100894
rect 207266 100338 207502 100574
rect 207586 100338 207822 100574
rect 207266 64658 207502 64894
rect 207586 64658 207822 64894
rect 207266 64338 207502 64574
rect 207586 64338 207822 64574
rect 207266 28658 207502 28894
rect 207586 28658 207822 28894
rect 207266 28338 207502 28574
rect 207586 28338 207822 28574
rect 207266 -5382 207502 -5146
rect 207586 -5382 207822 -5146
rect 207266 -5702 207502 -5466
rect 207586 -5702 207822 -5466
rect 228986 710362 229222 710598
rect 229306 710362 229542 710598
rect 228986 710042 229222 710278
rect 229306 710042 229542 710278
rect 225266 708442 225502 708678
rect 225586 708442 225822 708678
rect 225266 708122 225502 708358
rect 225586 708122 225822 708358
rect 221546 706522 221782 706758
rect 221866 706522 222102 706758
rect 221546 706202 221782 706438
rect 221866 706202 222102 706438
rect 210986 680378 211222 680614
rect 211306 680378 211542 680614
rect 210986 680058 211222 680294
rect 211306 680058 211542 680294
rect 210986 644378 211222 644614
rect 211306 644378 211542 644614
rect 210986 644058 211222 644294
rect 211306 644058 211542 644294
rect 210986 608378 211222 608614
rect 211306 608378 211542 608614
rect 210986 608058 211222 608294
rect 211306 608058 211542 608294
rect 210986 572378 211222 572614
rect 211306 572378 211542 572614
rect 210986 572058 211222 572294
rect 211306 572058 211542 572294
rect 210986 536378 211222 536614
rect 211306 536378 211542 536614
rect 210986 536058 211222 536294
rect 211306 536058 211542 536294
rect 210986 500378 211222 500614
rect 211306 500378 211542 500614
rect 210986 500058 211222 500294
rect 211306 500058 211542 500294
rect 210986 464378 211222 464614
rect 211306 464378 211542 464614
rect 210986 464058 211222 464294
rect 211306 464058 211542 464294
rect 210986 428378 211222 428614
rect 211306 428378 211542 428614
rect 210986 428058 211222 428294
rect 211306 428058 211542 428294
rect 210986 392378 211222 392614
rect 211306 392378 211542 392614
rect 210986 392058 211222 392294
rect 211306 392058 211542 392294
rect 210986 356378 211222 356614
rect 211306 356378 211542 356614
rect 210986 356058 211222 356294
rect 211306 356058 211542 356294
rect 210986 320378 211222 320614
rect 211306 320378 211542 320614
rect 210986 320058 211222 320294
rect 211306 320058 211542 320294
rect 210986 284378 211222 284614
rect 211306 284378 211542 284614
rect 210986 284058 211222 284294
rect 211306 284058 211542 284294
rect 210986 248378 211222 248614
rect 211306 248378 211542 248614
rect 210986 248058 211222 248294
rect 211306 248058 211542 248294
rect 210986 212378 211222 212614
rect 211306 212378 211542 212614
rect 210986 212058 211222 212294
rect 211306 212058 211542 212294
rect 210986 176378 211222 176614
rect 211306 176378 211542 176614
rect 210986 176058 211222 176294
rect 211306 176058 211542 176294
rect 210986 140378 211222 140614
rect 211306 140378 211542 140614
rect 210986 140058 211222 140294
rect 211306 140058 211542 140294
rect 210986 104378 211222 104614
rect 211306 104378 211542 104614
rect 210986 104058 211222 104294
rect 211306 104058 211542 104294
rect 210986 68378 211222 68614
rect 211306 68378 211542 68614
rect 210986 68058 211222 68294
rect 211306 68058 211542 68294
rect 210986 32378 211222 32614
rect 211306 32378 211542 32614
rect 210986 32058 211222 32294
rect 211306 32058 211542 32294
rect 192986 -6342 193222 -6106
rect 193306 -6342 193542 -6106
rect 192986 -6662 193222 -6426
rect 193306 -6662 193542 -6426
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 217826 543218 218062 543454
rect 218146 543218 218382 543454
rect 217826 542898 218062 543134
rect 218146 542898 218382 543134
rect 217826 507218 218062 507454
rect 218146 507218 218382 507454
rect 217826 506898 218062 507134
rect 218146 506898 218382 507134
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 217826 435218 218062 435454
rect 218146 435218 218382 435454
rect 217826 434898 218062 435134
rect 218146 434898 218382 435134
rect 217826 399218 218062 399454
rect 218146 399218 218382 399454
rect 217826 398898 218062 399134
rect 218146 398898 218382 399134
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 217826 327218 218062 327454
rect 218146 327218 218382 327454
rect 217826 326898 218062 327134
rect 218146 326898 218382 327134
rect 217826 291218 218062 291454
rect 218146 291218 218382 291454
rect 217826 290898 218062 291134
rect 218146 290898 218382 291134
rect 217826 255218 218062 255454
rect 218146 255218 218382 255454
rect 217826 254898 218062 255134
rect 218146 254898 218382 255134
rect 217826 219218 218062 219454
rect 218146 219218 218382 219454
rect 217826 218898 218062 219134
rect 218146 218898 218382 219134
rect 217826 183218 218062 183454
rect 218146 183218 218382 183454
rect 217826 182898 218062 183134
rect 218146 182898 218382 183134
rect 217826 147218 218062 147454
rect 218146 147218 218382 147454
rect 217826 146898 218062 147134
rect 218146 146898 218382 147134
rect 217826 111218 218062 111454
rect 218146 111218 218382 111454
rect 217826 110898 218062 111134
rect 218146 110898 218382 111134
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 221546 690938 221782 691174
rect 221866 690938 222102 691174
rect 221546 690618 221782 690854
rect 221866 690618 222102 690854
rect 221546 654938 221782 655174
rect 221866 654938 222102 655174
rect 221546 654618 221782 654854
rect 221866 654618 222102 654854
rect 221546 618938 221782 619174
rect 221866 618938 222102 619174
rect 221546 618618 221782 618854
rect 221866 618618 222102 618854
rect 221546 582938 221782 583174
rect 221866 582938 222102 583174
rect 221546 582618 221782 582854
rect 221866 582618 222102 582854
rect 221546 546938 221782 547174
rect 221866 546938 222102 547174
rect 221546 546618 221782 546854
rect 221866 546618 222102 546854
rect 221546 510938 221782 511174
rect 221866 510938 222102 511174
rect 221546 510618 221782 510854
rect 221866 510618 222102 510854
rect 221546 474938 221782 475174
rect 221866 474938 222102 475174
rect 221546 474618 221782 474854
rect 221866 474618 222102 474854
rect 221546 438938 221782 439174
rect 221866 438938 222102 439174
rect 221546 438618 221782 438854
rect 221866 438618 222102 438854
rect 221546 402938 221782 403174
rect 221866 402938 222102 403174
rect 221546 402618 221782 402854
rect 221866 402618 222102 402854
rect 221546 366938 221782 367174
rect 221866 366938 222102 367174
rect 221546 366618 221782 366854
rect 221866 366618 222102 366854
rect 221546 330938 221782 331174
rect 221866 330938 222102 331174
rect 221546 330618 221782 330854
rect 221866 330618 222102 330854
rect 221546 294938 221782 295174
rect 221866 294938 222102 295174
rect 221546 294618 221782 294854
rect 221866 294618 222102 294854
rect 221546 258938 221782 259174
rect 221866 258938 222102 259174
rect 221546 258618 221782 258854
rect 221866 258618 222102 258854
rect 221546 222938 221782 223174
rect 221866 222938 222102 223174
rect 221546 222618 221782 222854
rect 221866 222618 222102 222854
rect 221546 186938 221782 187174
rect 221866 186938 222102 187174
rect 221546 186618 221782 186854
rect 221866 186618 222102 186854
rect 221546 150938 221782 151174
rect 221866 150938 222102 151174
rect 221546 150618 221782 150854
rect 221866 150618 222102 150854
rect 221546 114938 221782 115174
rect 221866 114938 222102 115174
rect 221546 114618 221782 114854
rect 221866 114618 222102 114854
rect 221546 78938 221782 79174
rect 221866 78938 222102 79174
rect 221546 78618 221782 78854
rect 221866 78618 222102 78854
rect 221546 42938 221782 43174
rect 221866 42938 222102 43174
rect 221546 42618 221782 42854
rect 221866 42618 222102 42854
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 221546 -2502 221782 -2266
rect 221866 -2502 222102 -2266
rect 221546 -2822 221782 -2586
rect 221866 -2822 222102 -2586
rect 225266 694658 225502 694894
rect 225586 694658 225822 694894
rect 225266 694338 225502 694574
rect 225586 694338 225822 694574
rect 225266 658658 225502 658894
rect 225586 658658 225822 658894
rect 225266 658338 225502 658574
rect 225586 658338 225822 658574
rect 225266 622658 225502 622894
rect 225586 622658 225822 622894
rect 225266 622338 225502 622574
rect 225586 622338 225822 622574
rect 225266 586658 225502 586894
rect 225586 586658 225822 586894
rect 225266 586338 225502 586574
rect 225586 586338 225822 586574
rect 225266 550658 225502 550894
rect 225586 550658 225822 550894
rect 225266 550338 225502 550574
rect 225586 550338 225822 550574
rect 225266 514658 225502 514894
rect 225586 514658 225822 514894
rect 225266 514338 225502 514574
rect 225586 514338 225822 514574
rect 225266 478658 225502 478894
rect 225586 478658 225822 478894
rect 225266 478338 225502 478574
rect 225586 478338 225822 478574
rect 225266 442658 225502 442894
rect 225586 442658 225822 442894
rect 225266 442338 225502 442574
rect 225586 442338 225822 442574
rect 225266 406658 225502 406894
rect 225586 406658 225822 406894
rect 225266 406338 225502 406574
rect 225586 406338 225822 406574
rect 225266 370658 225502 370894
rect 225586 370658 225822 370894
rect 225266 370338 225502 370574
rect 225586 370338 225822 370574
rect 225266 334658 225502 334894
rect 225586 334658 225822 334894
rect 225266 334338 225502 334574
rect 225586 334338 225822 334574
rect 225266 298658 225502 298894
rect 225586 298658 225822 298894
rect 225266 298338 225502 298574
rect 225586 298338 225822 298574
rect 225266 262658 225502 262894
rect 225586 262658 225822 262894
rect 225266 262338 225502 262574
rect 225586 262338 225822 262574
rect 225266 226658 225502 226894
rect 225586 226658 225822 226894
rect 225266 226338 225502 226574
rect 225586 226338 225822 226574
rect 225266 190658 225502 190894
rect 225586 190658 225822 190894
rect 225266 190338 225502 190574
rect 225586 190338 225822 190574
rect 225266 154658 225502 154894
rect 225586 154658 225822 154894
rect 225266 154338 225502 154574
rect 225586 154338 225822 154574
rect 225266 118658 225502 118894
rect 225586 118658 225822 118894
rect 225266 118338 225502 118574
rect 225586 118338 225822 118574
rect 225266 82658 225502 82894
rect 225586 82658 225822 82894
rect 225266 82338 225502 82574
rect 225586 82338 225822 82574
rect 225266 46658 225502 46894
rect 225586 46658 225822 46894
rect 225266 46338 225502 46574
rect 225586 46338 225822 46574
rect 225266 10658 225502 10894
rect 225586 10658 225822 10894
rect 225266 10338 225502 10574
rect 225586 10338 225822 10574
rect 225266 -4422 225502 -4186
rect 225586 -4422 225822 -4186
rect 225266 -4742 225502 -4506
rect 225586 -4742 225822 -4506
rect 246986 711322 247222 711558
rect 247306 711322 247542 711558
rect 246986 711002 247222 711238
rect 247306 711002 247542 711238
rect 243266 709402 243502 709638
rect 243586 709402 243822 709638
rect 243266 709082 243502 709318
rect 243586 709082 243822 709318
rect 239546 707482 239782 707718
rect 239866 707482 240102 707718
rect 239546 707162 239782 707398
rect 239866 707162 240102 707398
rect 228986 698378 229222 698614
rect 229306 698378 229542 698614
rect 228986 698058 229222 698294
rect 229306 698058 229542 698294
rect 228986 662378 229222 662614
rect 229306 662378 229542 662614
rect 228986 662058 229222 662294
rect 229306 662058 229542 662294
rect 228986 626378 229222 626614
rect 229306 626378 229542 626614
rect 228986 626058 229222 626294
rect 229306 626058 229542 626294
rect 228986 590378 229222 590614
rect 229306 590378 229542 590614
rect 228986 590058 229222 590294
rect 229306 590058 229542 590294
rect 228986 554378 229222 554614
rect 229306 554378 229542 554614
rect 228986 554058 229222 554294
rect 229306 554058 229542 554294
rect 228986 518378 229222 518614
rect 229306 518378 229542 518614
rect 228986 518058 229222 518294
rect 229306 518058 229542 518294
rect 228986 482378 229222 482614
rect 229306 482378 229542 482614
rect 228986 482058 229222 482294
rect 229306 482058 229542 482294
rect 228986 446378 229222 446614
rect 229306 446378 229542 446614
rect 228986 446058 229222 446294
rect 229306 446058 229542 446294
rect 228986 410378 229222 410614
rect 229306 410378 229542 410614
rect 228986 410058 229222 410294
rect 229306 410058 229542 410294
rect 228986 374378 229222 374614
rect 229306 374378 229542 374614
rect 228986 374058 229222 374294
rect 229306 374058 229542 374294
rect 235826 705562 236062 705798
rect 236146 705562 236382 705798
rect 235826 705242 236062 705478
rect 236146 705242 236382 705478
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 235826 561218 236062 561454
rect 236146 561218 236382 561454
rect 235826 560898 236062 561134
rect 236146 560898 236382 561134
rect 235826 525218 236062 525454
rect 236146 525218 236382 525454
rect 235826 524898 236062 525134
rect 236146 524898 236382 525134
rect 235826 489218 236062 489454
rect 236146 489218 236382 489454
rect 235826 488898 236062 489134
rect 236146 488898 236382 489134
rect 235826 453218 236062 453454
rect 236146 453218 236382 453454
rect 235826 452898 236062 453134
rect 236146 452898 236382 453134
rect 235826 417218 236062 417454
rect 236146 417218 236382 417454
rect 235826 416898 236062 417134
rect 236146 416898 236382 417134
rect 235826 381218 236062 381454
rect 236146 381218 236382 381454
rect 235826 380898 236062 381134
rect 236146 380898 236382 381134
rect 235826 345218 236062 345454
rect 236146 345218 236382 345454
rect 228986 338378 229222 338614
rect 229306 338378 229542 338614
rect 228986 338058 229222 338294
rect 229306 338058 229542 338294
rect 228986 302378 229222 302614
rect 229306 302378 229542 302614
rect 228986 302058 229222 302294
rect 229306 302058 229542 302294
rect 228986 266378 229222 266614
rect 229306 266378 229542 266614
rect 228986 266058 229222 266294
rect 229306 266058 229542 266294
rect 228986 230378 229222 230614
rect 229306 230378 229542 230614
rect 228986 230058 229222 230294
rect 229306 230058 229542 230294
rect 228986 194378 229222 194614
rect 229306 194378 229542 194614
rect 228986 194058 229222 194294
rect 229306 194058 229542 194294
rect 235826 344898 236062 345134
rect 236146 344898 236382 345134
rect 235826 309218 236062 309454
rect 236146 309218 236382 309454
rect 235826 308898 236062 309134
rect 236146 308898 236382 309134
rect 235826 273218 236062 273454
rect 236146 273218 236382 273454
rect 235826 272898 236062 273134
rect 236146 272898 236382 273134
rect 235826 237218 236062 237454
rect 236146 237218 236382 237454
rect 235826 236898 236062 237134
rect 236146 236898 236382 237134
rect 235826 201218 236062 201454
rect 236146 201218 236382 201454
rect 235826 200898 236062 201134
rect 236146 200898 236382 201134
rect 228986 158378 229222 158614
rect 229306 158378 229542 158614
rect 228986 158058 229222 158294
rect 229306 158058 229542 158294
rect 228986 122378 229222 122614
rect 229306 122378 229542 122614
rect 228986 122058 229222 122294
rect 229306 122058 229542 122294
rect 228986 86378 229222 86614
rect 229306 86378 229542 86614
rect 228986 86058 229222 86294
rect 229306 86058 229542 86294
rect 228986 50378 229222 50614
rect 229306 50378 229542 50614
rect 228986 50058 229222 50294
rect 229306 50058 229542 50294
rect 228986 14378 229222 14614
rect 229306 14378 229542 14614
rect 228986 14058 229222 14294
rect 229306 14058 229542 14294
rect 210986 -7302 211222 -7066
rect 211306 -7302 211542 -7066
rect 210986 -7622 211222 -7386
rect 211306 -7622 211542 -7386
rect 239546 672938 239782 673174
rect 239866 672938 240102 673174
rect 239546 672618 239782 672854
rect 239866 672618 240102 672854
rect 239546 636938 239782 637174
rect 239866 636938 240102 637174
rect 239546 636618 239782 636854
rect 239866 636618 240102 636854
rect 239546 600938 239782 601174
rect 239866 600938 240102 601174
rect 239546 600618 239782 600854
rect 239866 600618 240102 600854
rect 239546 564938 239782 565174
rect 239866 564938 240102 565174
rect 239546 564618 239782 564854
rect 239866 564618 240102 564854
rect 239546 528938 239782 529174
rect 239866 528938 240102 529174
rect 239546 528618 239782 528854
rect 239866 528618 240102 528854
rect 239546 492938 239782 493174
rect 239866 492938 240102 493174
rect 239546 492618 239782 492854
rect 239866 492618 240102 492854
rect 239546 456938 239782 457174
rect 239866 456938 240102 457174
rect 239546 456618 239782 456854
rect 239866 456618 240102 456854
rect 243266 676658 243502 676894
rect 243586 676658 243822 676894
rect 243266 676338 243502 676574
rect 243586 676338 243822 676574
rect 243266 640658 243502 640894
rect 243586 640658 243822 640894
rect 243266 640338 243502 640574
rect 243586 640338 243822 640574
rect 243266 604658 243502 604894
rect 243586 604658 243822 604894
rect 243266 604338 243502 604574
rect 243586 604338 243822 604574
rect 243266 568658 243502 568894
rect 243586 568658 243822 568894
rect 243266 568338 243502 568574
rect 243586 568338 243822 568574
rect 243266 532658 243502 532894
rect 243586 532658 243822 532894
rect 243266 532338 243502 532574
rect 243586 532338 243822 532574
rect 243266 496658 243502 496894
rect 243586 496658 243822 496894
rect 243266 496338 243502 496574
rect 243586 496338 243822 496574
rect 243266 460658 243502 460894
rect 243586 460658 243822 460894
rect 243266 460338 243502 460574
rect 243586 460338 243822 460574
rect 264986 710362 265222 710598
rect 265306 710362 265542 710598
rect 264986 710042 265222 710278
rect 265306 710042 265542 710278
rect 261266 708442 261502 708678
rect 261586 708442 261822 708678
rect 261266 708122 261502 708358
rect 261586 708122 261822 708358
rect 257546 706522 257782 706758
rect 257866 706522 258102 706758
rect 257546 706202 257782 706438
rect 257866 706202 258102 706438
rect 246986 680378 247222 680614
rect 247306 680378 247542 680614
rect 246986 680058 247222 680294
rect 247306 680058 247542 680294
rect 246986 644378 247222 644614
rect 247306 644378 247542 644614
rect 246986 644058 247222 644294
rect 247306 644058 247542 644294
rect 246986 608378 247222 608614
rect 247306 608378 247542 608614
rect 246986 608058 247222 608294
rect 247306 608058 247542 608294
rect 246986 572378 247222 572614
rect 247306 572378 247542 572614
rect 246986 572058 247222 572294
rect 247306 572058 247542 572294
rect 246986 536378 247222 536614
rect 247306 536378 247542 536614
rect 246986 536058 247222 536294
rect 247306 536058 247542 536294
rect 246986 500378 247222 500614
rect 247306 500378 247542 500614
rect 246986 500058 247222 500294
rect 247306 500058 247542 500294
rect 246986 464378 247222 464614
rect 247306 464378 247542 464614
rect 246986 464058 247222 464294
rect 247306 464058 247542 464294
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 253826 543218 254062 543454
rect 254146 543218 254382 543454
rect 253826 542898 254062 543134
rect 254146 542898 254382 543134
rect 253826 507218 254062 507454
rect 254146 507218 254382 507454
rect 253826 506898 254062 507134
rect 254146 506898 254382 507134
rect 253826 471218 254062 471454
rect 254146 471218 254382 471454
rect 253826 470898 254062 471134
rect 254146 470898 254382 471134
rect 257546 690938 257782 691174
rect 257866 690938 258102 691174
rect 257546 690618 257782 690854
rect 257866 690618 258102 690854
rect 257546 654938 257782 655174
rect 257866 654938 258102 655174
rect 257546 654618 257782 654854
rect 257866 654618 258102 654854
rect 257546 618938 257782 619174
rect 257866 618938 258102 619174
rect 257546 618618 257782 618854
rect 257866 618618 258102 618854
rect 257546 582938 257782 583174
rect 257866 582938 258102 583174
rect 257546 582618 257782 582854
rect 257866 582618 258102 582854
rect 257546 546938 257782 547174
rect 257866 546938 258102 547174
rect 257546 546618 257782 546854
rect 257866 546618 258102 546854
rect 257546 510938 257782 511174
rect 257866 510938 258102 511174
rect 257546 510618 257782 510854
rect 257866 510618 258102 510854
rect 257546 474938 257782 475174
rect 257866 474938 258102 475174
rect 257546 474618 257782 474854
rect 257866 474618 258102 474854
rect 261266 694658 261502 694894
rect 261586 694658 261822 694894
rect 261266 694338 261502 694574
rect 261586 694338 261822 694574
rect 261266 658658 261502 658894
rect 261586 658658 261822 658894
rect 261266 658338 261502 658574
rect 261586 658338 261822 658574
rect 261266 622658 261502 622894
rect 261586 622658 261822 622894
rect 261266 622338 261502 622574
rect 261586 622338 261822 622574
rect 261266 586658 261502 586894
rect 261586 586658 261822 586894
rect 261266 586338 261502 586574
rect 261586 586338 261822 586574
rect 261266 550658 261502 550894
rect 261586 550658 261822 550894
rect 261266 550338 261502 550574
rect 261586 550338 261822 550574
rect 261266 514658 261502 514894
rect 261586 514658 261822 514894
rect 261266 514338 261502 514574
rect 261586 514338 261822 514574
rect 261266 478658 261502 478894
rect 261586 478658 261822 478894
rect 261266 478338 261502 478574
rect 261586 478338 261822 478574
rect 261266 442658 261502 442894
rect 261586 442658 261822 442894
rect 261266 442338 261502 442574
rect 261586 442338 261822 442574
rect 282986 711322 283222 711558
rect 283306 711322 283542 711558
rect 282986 711002 283222 711238
rect 283306 711002 283542 711238
rect 279266 709402 279502 709638
rect 279586 709402 279822 709638
rect 279266 709082 279502 709318
rect 279586 709082 279822 709318
rect 275546 707482 275782 707718
rect 275866 707482 276102 707718
rect 275546 707162 275782 707398
rect 275866 707162 276102 707398
rect 264986 698378 265222 698614
rect 265306 698378 265542 698614
rect 264986 698058 265222 698294
rect 265306 698058 265542 698294
rect 264986 662378 265222 662614
rect 265306 662378 265542 662614
rect 264986 662058 265222 662294
rect 265306 662058 265542 662294
rect 264986 626378 265222 626614
rect 265306 626378 265542 626614
rect 264986 626058 265222 626294
rect 265306 626058 265542 626294
rect 264986 590378 265222 590614
rect 265306 590378 265542 590614
rect 264986 590058 265222 590294
rect 265306 590058 265542 590294
rect 264986 554378 265222 554614
rect 265306 554378 265542 554614
rect 264986 554058 265222 554294
rect 265306 554058 265542 554294
rect 264986 518378 265222 518614
rect 265306 518378 265542 518614
rect 264986 518058 265222 518294
rect 265306 518058 265542 518294
rect 264986 482378 265222 482614
rect 265306 482378 265542 482614
rect 264986 482058 265222 482294
rect 265306 482058 265542 482294
rect 264986 446378 265222 446614
rect 265306 446378 265542 446614
rect 264986 446058 265222 446294
rect 265306 446058 265542 446294
rect 271826 705562 272062 705798
rect 272146 705562 272382 705798
rect 271826 705242 272062 705478
rect 272146 705242 272382 705478
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 271826 561218 272062 561454
rect 272146 561218 272382 561454
rect 271826 560898 272062 561134
rect 272146 560898 272382 561134
rect 271826 525218 272062 525454
rect 272146 525218 272382 525454
rect 271826 524898 272062 525134
rect 272146 524898 272382 525134
rect 271826 489218 272062 489454
rect 272146 489218 272382 489454
rect 271826 488898 272062 489134
rect 272146 488898 272382 489134
rect 271826 453218 272062 453454
rect 272146 453218 272382 453454
rect 271826 452898 272062 453134
rect 272146 452898 272382 453134
rect 275546 672938 275782 673174
rect 275866 672938 276102 673174
rect 275546 672618 275782 672854
rect 275866 672618 276102 672854
rect 275546 636938 275782 637174
rect 275866 636938 276102 637174
rect 275546 636618 275782 636854
rect 275866 636618 276102 636854
rect 275546 600938 275782 601174
rect 275866 600938 276102 601174
rect 275546 600618 275782 600854
rect 275866 600618 276102 600854
rect 275546 564938 275782 565174
rect 275866 564938 276102 565174
rect 275546 564618 275782 564854
rect 275866 564618 276102 564854
rect 275546 528938 275782 529174
rect 275866 528938 276102 529174
rect 275546 528618 275782 528854
rect 275866 528618 276102 528854
rect 275546 492938 275782 493174
rect 275866 492938 276102 493174
rect 275546 492618 275782 492854
rect 275866 492618 276102 492854
rect 275546 456938 275782 457174
rect 275866 456938 276102 457174
rect 275546 456618 275782 456854
rect 275866 456618 276102 456854
rect 279266 676658 279502 676894
rect 279586 676658 279822 676894
rect 279266 676338 279502 676574
rect 279586 676338 279822 676574
rect 279266 640658 279502 640894
rect 279586 640658 279822 640894
rect 279266 640338 279502 640574
rect 279586 640338 279822 640574
rect 279266 604658 279502 604894
rect 279586 604658 279822 604894
rect 279266 604338 279502 604574
rect 279586 604338 279822 604574
rect 279266 568658 279502 568894
rect 279586 568658 279822 568894
rect 279266 568338 279502 568574
rect 279586 568338 279822 568574
rect 279266 532658 279502 532894
rect 279586 532658 279822 532894
rect 279266 532338 279502 532574
rect 279586 532338 279822 532574
rect 279266 496658 279502 496894
rect 279586 496658 279822 496894
rect 279266 496338 279502 496574
rect 279586 496338 279822 496574
rect 279266 460658 279502 460894
rect 279586 460658 279822 460894
rect 279266 460338 279502 460574
rect 279586 460338 279822 460574
rect 300986 710362 301222 710598
rect 301306 710362 301542 710598
rect 300986 710042 301222 710278
rect 301306 710042 301542 710278
rect 297266 708442 297502 708678
rect 297586 708442 297822 708678
rect 297266 708122 297502 708358
rect 297586 708122 297822 708358
rect 293546 706522 293782 706758
rect 293866 706522 294102 706758
rect 293546 706202 293782 706438
rect 293866 706202 294102 706438
rect 282986 680378 283222 680614
rect 283306 680378 283542 680614
rect 282986 680058 283222 680294
rect 283306 680058 283542 680294
rect 282986 644378 283222 644614
rect 283306 644378 283542 644614
rect 282986 644058 283222 644294
rect 283306 644058 283542 644294
rect 282986 608378 283222 608614
rect 283306 608378 283542 608614
rect 282986 608058 283222 608294
rect 283306 608058 283542 608294
rect 282986 572378 283222 572614
rect 283306 572378 283542 572614
rect 282986 572058 283222 572294
rect 283306 572058 283542 572294
rect 282986 536378 283222 536614
rect 283306 536378 283542 536614
rect 282986 536058 283222 536294
rect 283306 536058 283542 536294
rect 282986 500378 283222 500614
rect 283306 500378 283542 500614
rect 282986 500058 283222 500294
rect 283306 500058 283542 500294
rect 282986 464378 283222 464614
rect 283306 464378 283542 464614
rect 282986 464058 283222 464294
rect 283306 464058 283542 464294
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 289826 507218 290062 507454
rect 290146 507218 290382 507454
rect 289826 506898 290062 507134
rect 290146 506898 290382 507134
rect 289826 471218 290062 471454
rect 290146 471218 290382 471454
rect 289826 470898 290062 471134
rect 290146 470898 290382 471134
rect 293546 690938 293782 691174
rect 293866 690938 294102 691174
rect 293546 690618 293782 690854
rect 293866 690618 294102 690854
rect 293546 654938 293782 655174
rect 293866 654938 294102 655174
rect 293546 654618 293782 654854
rect 293866 654618 294102 654854
rect 293546 618938 293782 619174
rect 293866 618938 294102 619174
rect 293546 618618 293782 618854
rect 293866 618618 294102 618854
rect 293546 582938 293782 583174
rect 293866 582938 294102 583174
rect 293546 582618 293782 582854
rect 293866 582618 294102 582854
rect 293546 546938 293782 547174
rect 293866 546938 294102 547174
rect 293546 546618 293782 546854
rect 293866 546618 294102 546854
rect 293546 510938 293782 511174
rect 293866 510938 294102 511174
rect 293546 510618 293782 510854
rect 293866 510618 294102 510854
rect 293546 474938 293782 475174
rect 293866 474938 294102 475174
rect 293546 474618 293782 474854
rect 293866 474618 294102 474854
rect 297266 694658 297502 694894
rect 297586 694658 297822 694894
rect 297266 694338 297502 694574
rect 297586 694338 297822 694574
rect 297266 658658 297502 658894
rect 297586 658658 297822 658894
rect 297266 658338 297502 658574
rect 297586 658338 297822 658574
rect 297266 622658 297502 622894
rect 297586 622658 297822 622894
rect 297266 622338 297502 622574
rect 297586 622338 297822 622574
rect 297266 586658 297502 586894
rect 297586 586658 297822 586894
rect 297266 586338 297502 586574
rect 297586 586338 297822 586574
rect 297266 550658 297502 550894
rect 297586 550658 297822 550894
rect 297266 550338 297502 550574
rect 297586 550338 297822 550574
rect 297266 514658 297502 514894
rect 297586 514658 297822 514894
rect 297266 514338 297502 514574
rect 297586 514338 297822 514574
rect 297266 478658 297502 478894
rect 297586 478658 297822 478894
rect 297266 478338 297502 478574
rect 297586 478338 297822 478574
rect 297266 442658 297502 442894
rect 297586 442658 297822 442894
rect 297266 442338 297502 442574
rect 297586 442338 297822 442574
rect 318986 711322 319222 711558
rect 319306 711322 319542 711558
rect 318986 711002 319222 711238
rect 319306 711002 319542 711238
rect 315266 709402 315502 709638
rect 315586 709402 315822 709638
rect 315266 709082 315502 709318
rect 315586 709082 315822 709318
rect 311546 707482 311782 707718
rect 311866 707482 312102 707718
rect 311546 707162 311782 707398
rect 311866 707162 312102 707398
rect 300986 698378 301222 698614
rect 301306 698378 301542 698614
rect 300986 698058 301222 698294
rect 301306 698058 301542 698294
rect 300986 662378 301222 662614
rect 301306 662378 301542 662614
rect 300986 662058 301222 662294
rect 301306 662058 301542 662294
rect 300986 626378 301222 626614
rect 301306 626378 301542 626614
rect 300986 626058 301222 626294
rect 301306 626058 301542 626294
rect 300986 590378 301222 590614
rect 301306 590378 301542 590614
rect 300986 590058 301222 590294
rect 301306 590058 301542 590294
rect 300986 554378 301222 554614
rect 301306 554378 301542 554614
rect 300986 554058 301222 554294
rect 301306 554058 301542 554294
rect 300986 518378 301222 518614
rect 301306 518378 301542 518614
rect 300986 518058 301222 518294
rect 301306 518058 301542 518294
rect 300986 482378 301222 482614
rect 301306 482378 301542 482614
rect 300986 482058 301222 482294
rect 301306 482058 301542 482294
rect 300986 446378 301222 446614
rect 301306 446378 301542 446614
rect 300986 446058 301222 446294
rect 301306 446058 301542 446294
rect 307826 705562 308062 705798
rect 308146 705562 308382 705798
rect 307826 705242 308062 705478
rect 308146 705242 308382 705478
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 307826 561218 308062 561454
rect 308146 561218 308382 561454
rect 307826 560898 308062 561134
rect 308146 560898 308382 561134
rect 307826 525218 308062 525454
rect 308146 525218 308382 525454
rect 307826 524898 308062 525134
rect 308146 524898 308382 525134
rect 307826 489218 308062 489454
rect 308146 489218 308382 489454
rect 307826 488898 308062 489134
rect 308146 488898 308382 489134
rect 307826 453218 308062 453454
rect 308146 453218 308382 453454
rect 307826 452898 308062 453134
rect 308146 452898 308382 453134
rect 311546 672938 311782 673174
rect 311866 672938 312102 673174
rect 311546 672618 311782 672854
rect 311866 672618 312102 672854
rect 311546 636938 311782 637174
rect 311866 636938 312102 637174
rect 311546 636618 311782 636854
rect 311866 636618 312102 636854
rect 311546 600938 311782 601174
rect 311866 600938 312102 601174
rect 311546 600618 311782 600854
rect 311866 600618 312102 600854
rect 311546 564938 311782 565174
rect 311866 564938 312102 565174
rect 311546 564618 311782 564854
rect 311866 564618 312102 564854
rect 311546 528938 311782 529174
rect 311866 528938 312102 529174
rect 311546 528618 311782 528854
rect 311866 528618 312102 528854
rect 311546 492938 311782 493174
rect 311866 492938 312102 493174
rect 311546 492618 311782 492854
rect 311866 492618 312102 492854
rect 311546 456938 311782 457174
rect 311866 456938 312102 457174
rect 311546 456618 311782 456854
rect 311866 456618 312102 456854
rect 315266 676658 315502 676894
rect 315586 676658 315822 676894
rect 315266 676338 315502 676574
rect 315586 676338 315822 676574
rect 315266 640658 315502 640894
rect 315586 640658 315822 640894
rect 315266 640338 315502 640574
rect 315586 640338 315822 640574
rect 315266 604658 315502 604894
rect 315586 604658 315822 604894
rect 315266 604338 315502 604574
rect 315586 604338 315822 604574
rect 315266 568658 315502 568894
rect 315586 568658 315822 568894
rect 315266 568338 315502 568574
rect 315586 568338 315822 568574
rect 315266 532658 315502 532894
rect 315586 532658 315822 532894
rect 315266 532338 315502 532574
rect 315586 532338 315822 532574
rect 315266 496658 315502 496894
rect 315586 496658 315822 496894
rect 315266 496338 315502 496574
rect 315586 496338 315822 496574
rect 315266 460658 315502 460894
rect 315586 460658 315822 460894
rect 315266 460338 315502 460574
rect 315586 460338 315822 460574
rect 336986 710362 337222 710598
rect 337306 710362 337542 710598
rect 336986 710042 337222 710278
rect 337306 710042 337542 710278
rect 333266 708442 333502 708678
rect 333586 708442 333822 708678
rect 333266 708122 333502 708358
rect 333586 708122 333822 708358
rect 329546 706522 329782 706758
rect 329866 706522 330102 706758
rect 329546 706202 329782 706438
rect 329866 706202 330102 706438
rect 318986 680378 319222 680614
rect 319306 680378 319542 680614
rect 318986 680058 319222 680294
rect 319306 680058 319542 680294
rect 318986 644378 319222 644614
rect 319306 644378 319542 644614
rect 318986 644058 319222 644294
rect 319306 644058 319542 644294
rect 318986 608378 319222 608614
rect 319306 608378 319542 608614
rect 318986 608058 319222 608294
rect 319306 608058 319542 608294
rect 318986 572378 319222 572614
rect 319306 572378 319542 572614
rect 318986 572058 319222 572294
rect 319306 572058 319542 572294
rect 318986 536378 319222 536614
rect 319306 536378 319542 536614
rect 318986 536058 319222 536294
rect 319306 536058 319542 536294
rect 318986 500378 319222 500614
rect 319306 500378 319542 500614
rect 318986 500058 319222 500294
rect 319306 500058 319542 500294
rect 318986 464378 319222 464614
rect 319306 464378 319542 464614
rect 318986 464058 319222 464294
rect 319306 464058 319542 464294
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 325826 543218 326062 543454
rect 326146 543218 326382 543454
rect 325826 542898 326062 543134
rect 326146 542898 326382 543134
rect 325826 507218 326062 507454
rect 326146 507218 326382 507454
rect 325826 506898 326062 507134
rect 326146 506898 326382 507134
rect 325826 471218 326062 471454
rect 326146 471218 326382 471454
rect 325826 470898 326062 471134
rect 326146 470898 326382 471134
rect 329546 690938 329782 691174
rect 329866 690938 330102 691174
rect 329546 690618 329782 690854
rect 329866 690618 330102 690854
rect 329546 654938 329782 655174
rect 329866 654938 330102 655174
rect 329546 654618 329782 654854
rect 329866 654618 330102 654854
rect 329546 618938 329782 619174
rect 329866 618938 330102 619174
rect 329546 618618 329782 618854
rect 329866 618618 330102 618854
rect 329546 582938 329782 583174
rect 329866 582938 330102 583174
rect 329546 582618 329782 582854
rect 329866 582618 330102 582854
rect 329546 546938 329782 547174
rect 329866 546938 330102 547174
rect 329546 546618 329782 546854
rect 329866 546618 330102 546854
rect 329546 510938 329782 511174
rect 329866 510938 330102 511174
rect 329546 510618 329782 510854
rect 329866 510618 330102 510854
rect 329546 474938 329782 475174
rect 329866 474938 330102 475174
rect 329546 474618 329782 474854
rect 329866 474618 330102 474854
rect 333266 694658 333502 694894
rect 333586 694658 333822 694894
rect 333266 694338 333502 694574
rect 333586 694338 333822 694574
rect 333266 658658 333502 658894
rect 333586 658658 333822 658894
rect 333266 658338 333502 658574
rect 333586 658338 333822 658574
rect 333266 622658 333502 622894
rect 333586 622658 333822 622894
rect 333266 622338 333502 622574
rect 333586 622338 333822 622574
rect 333266 586658 333502 586894
rect 333586 586658 333822 586894
rect 333266 586338 333502 586574
rect 333586 586338 333822 586574
rect 333266 550658 333502 550894
rect 333586 550658 333822 550894
rect 333266 550338 333502 550574
rect 333586 550338 333822 550574
rect 333266 514658 333502 514894
rect 333586 514658 333822 514894
rect 333266 514338 333502 514574
rect 333586 514338 333822 514574
rect 333266 478658 333502 478894
rect 333586 478658 333822 478894
rect 333266 478338 333502 478574
rect 333586 478338 333822 478574
rect 333266 442658 333502 442894
rect 333586 442658 333822 442894
rect 333266 442338 333502 442574
rect 333586 442338 333822 442574
rect 354986 711322 355222 711558
rect 355306 711322 355542 711558
rect 354986 711002 355222 711238
rect 355306 711002 355542 711238
rect 351266 709402 351502 709638
rect 351586 709402 351822 709638
rect 351266 709082 351502 709318
rect 351586 709082 351822 709318
rect 347546 707482 347782 707718
rect 347866 707482 348102 707718
rect 347546 707162 347782 707398
rect 347866 707162 348102 707398
rect 336986 698378 337222 698614
rect 337306 698378 337542 698614
rect 336986 698058 337222 698294
rect 337306 698058 337542 698294
rect 336986 662378 337222 662614
rect 337306 662378 337542 662614
rect 336986 662058 337222 662294
rect 337306 662058 337542 662294
rect 336986 626378 337222 626614
rect 337306 626378 337542 626614
rect 336986 626058 337222 626294
rect 337306 626058 337542 626294
rect 336986 590378 337222 590614
rect 337306 590378 337542 590614
rect 336986 590058 337222 590294
rect 337306 590058 337542 590294
rect 336986 554378 337222 554614
rect 337306 554378 337542 554614
rect 336986 554058 337222 554294
rect 337306 554058 337542 554294
rect 336986 518378 337222 518614
rect 337306 518378 337542 518614
rect 336986 518058 337222 518294
rect 337306 518058 337542 518294
rect 336986 482378 337222 482614
rect 337306 482378 337542 482614
rect 336986 482058 337222 482294
rect 337306 482058 337542 482294
rect 336986 446378 337222 446614
rect 337306 446378 337542 446614
rect 336986 446058 337222 446294
rect 337306 446058 337542 446294
rect 343826 705562 344062 705798
rect 344146 705562 344382 705798
rect 343826 705242 344062 705478
rect 344146 705242 344382 705478
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 343826 561218 344062 561454
rect 344146 561218 344382 561454
rect 343826 560898 344062 561134
rect 344146 560898 344382 561134
rect 343826 525218 344062 525454
rect 344146 525218 344382 525454
rect 343826 524898 344062 525134
rect 344146 524898 344382 525134
rect 343826 489218 344062 489454
rect 344146 489218 344382 489454
rect 343826 488898 344062 489134
rect 344146 488898 344382 489134
rect 343826 453218 344062 453454
rect 344146 453218 344382 453454
rect 343826 452898 344062 453134
rect 344146 452898 344382 453134
rect 347546 672938 347782 673174
rect 347866 672938 348102 673174
rect 347546 672618 347782 672854
rect 347866 672618 348102 672854
rect 347546 636938 347782 637174
rect 347866 636938 348102 637174
rect 347546 636618 347782 636854
rect 347866 636618 348102 636854
rect 347546 600938 347782 601174
rect 347866 600938 348102 601174
rect 347546 600618 347782 600854
rect 347866 600618 348102 600854
rect 347546 564938 347782 565174
rect 347866 564938 348102 565174
rect 347546 564618 347782 564854
rect 347866 564618 348102 564854
rect 347546 528938 347782 529174
rect 347866 528938 348102 529174
rect 347546 528618 347782 528854
rect 347866 528618 348102 528854
rect 347546 492938 347782 493174
rect 347866 492938 348102 493174
rect 347546 492618 347782 492854
rect 347866 492618 348102 492854
rect 347546 456938 347782 457174
rect 347866 456938 348102 457174
rect 347546 456618 347782 456854
rect 347866 456618 348102 456854
rect 351266 676658 351502 676894
rect 351586 676658 351822 676894
rect 351266 676338 351502 676574
rect 351586 676338 351822 676574
rect 351266 640658 351502 640894
rect 351586 640658 351822 640894
rect 351266 640338 351502 640574
rect 351586 640338 351822 640574
rect 351266 604658 351502 604894
rect 351586 604658 351822 604894
rect 351266 604338 351502 604574
rect 351586 604338 351822 604574
rect 351266 568658 351502 568894
rect 351586 568658 351822 568894
rect 351266 568338 351502 568574
rect 351586 568338 351822 568574
rect 351266 532658 351502 532894
rect 351586 532658 351822 532894
rect 351266 532338 351502 532574
rect 351586 532338 351822 532574
rect 351266 496658 351502 496894
rect 351586 496658 351822 496894
rect 351266 496338 351502 496574
rect 351586 496338 351822 496574
rect 351266 460658 351502 460894
rect 351586 460658 351822 460894
rect 351266 460338 351502 460574
rect 351586 460338 351822 460574
rect 372986 710362 373222 710598
rect 373306 710362 373542 710598
rect 372986 710042 373222 710278
rect 373306 710042 373542 710278
rect 369266 708442 369502 708678
rect 369586 708442 369822 708678
rect 369266 708122 369502 708358
rect 369586 708122 369822 708358
rect 365546 706522 365782 706758
rect 365866 706522 366102 706758
rect 365546 706202 365782 706438
rect 365866 706202 366102 706438
rect 354986 680378 355222 680614
rect 355306 680378 355542 680614
rect 354986 680058 355222 680294
rect 355306 680058 355542 680294
rect 354986 644378 355222 644614
rect 355306 644378 355542 644614
rect 354986 644058 355222 644294
rect 355306 644058 355542 644294
rect 354986 608378 355222 608614
rect 355306 608378 355542 608614
rect 354986 608058 355222 608294
rect 355306 608058 355542 608294
rect 354986 572378 355222 572614
rect 355306 572378 355542 572614
rect 354986 572058 355222 572294
rect 355306 572058 355542 572294
rect 354986 536378 355222 536614
rect 355306 536378 355542 536614
rect 354986 536058 355222 536294
rect 355306 536058 355542 536294
rect 354986 500378 355222 500614
rect 355306 500378 355542 500614
rect 354986 500058 355222 500294
rect 355306 500058 355542 500294
rect 354986 464378 355222 464614
rect 355306 464378 355542 464614
rect 354986 464058 355222 464294
rect 355306 464058 355542 464294
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 365546 690938 365782 691174
rect 365866 690938 366102 691174
rect 365546 690618 365782 690854
rect 365866 690618 366102 690854
rect 365546 654938 365782 655174
rect 365866 654938 366102 655174
rect 365546 654618 365782 654854
rect 365866 654618 366102 654854
rect 365546 618938 365782 619174
rect 365866 618938 366102 619174
rect 365546 618618 365782 618854
rect 365866 618618 366102 618854
rect 365546 582938 365782 583174
rect 365866 582938 366102 583174
rect 365546 582618 365782 582854
rect 365866 582618 366102 582854
rect 365546 546938 365782 547174
rect 365866 546938 366102 547174
rect 365546 546618 365782 546854
rect 365866 546618 366102 546854
rect 365546 510938 365782 511174
rect 365866 510938 366102 511174
rect 365546 510618 365782 510854
rect 365866 510618 366102 510854
rect 365546 474938 365782 475174
rect 365866 474938 366102 475174
rect 365546 474618 365782 474854
rect 365866 474618 366102 474854
rect 369266 694658 369502 694894
rect 369586 694658 369822 694894
rect 369266 694338 369502 694574
rect 369586 694338 369822 694574
rect 369266 658658 369502 658894
rect 369586 658658 369822 658894
rect 369266 658338 369502 658574
rect 369586 658338 369822 658574
rect 369266 622658 369502 622894
rect 369586 622658 369822 622894
rect 369266 622338 369502 622574
rect 369586 622338 369822 622574
rect 369266 586658 369502 586894
rect 369586 586658 369822 586894
rect 369266 586338 369502 586574
rect 369586 586338 369822 586574
rect 369266 550658 369502 550894
rect 369586 550658 369822 550894
rect 369266 550338 369502 550574
rect 369586 550338 369822 550574
rect 369266 514658 369502 514894
rect 369586 514658 369822 514894
rect 369266 514338 369502 514574
rect 369586 514338 369822 514574
rect 369266 478658 369502 478894
rect 369586 478658 369822 478894
rect 369266 478338 369502 478574
rect 369586 478338 369822 478574
rect 369266 442658 369502 442894
rect 369586 442658 369822 442894
rect 369266 442338 369502 442574
rect 369586 442338 369822 442574
rect 390986 711322 391222 711558
rect 391306 711322 391542 711558
rect 390986 711002 391222 711238
rect 391306 711002 391542 711238
rect 387266 709402 387502 709638
rect 387586 709402 387822 709638
rect 387266 709082 387502 709318
rect 387586 709082 387822 709318
rect 383546 707482 383782 707718
rect 383866 707482 384102 707718
rect 383546 707162 383782 707398
rect 383866 707162 384102 707398
rect 372986 698378 373222 698614
rect 373306 698378 373542 698614
rect 372986 698058 373222 698294
rect 373306 698058 373542 698294
rect 372986 662378 373222 662614
rect 373306 662378 373542 662614
rect 372986 662058 373222 662294
rect 373306 662058 373542 662294
rect 372986 626378 373222 626614
rect 373306 626378 373542 626614
rect 372986 626058 373222 626294
rect 373306 626058 373542 626294
rect 372986 590378 373222 590614
rect 373306 590378 373542 590614
rect 372986 590058 373222 590294
rect 373306 590058 373542 590294
rect 372986 554378 373222 554614
rect 373306 554378 373542 554614
rect 372986 554058 373222 554294
rect 373306 554058 373542 554294
rect 372986 518378 373222 518614
rect 373306 518378 373542 518614
rect 372986 518058 373222 518294
rect 373306 518058 373542 518294
rect 372986 482378 373222 482614
rect 373306 482378 373542 482614
rect 372986 482058 373222 482294
rect 373306 482058 373542 482294
rect 372986 446378 373222 446614
rect 373306 446378 373542 446614
rect 372986 446058 373222 446294
rect 373306 446058 373542 446294
rect 379826 705562 380062 705798
rect 380146 705562 380382 705798
rect 379826 705242 380062 705478
rect 380146 705242 380382 705478
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 379826 561218 380062 561454
rect 380146 561218 380382 561454
rect 379826 560898 380062 561134
rect 380146 560898 380382 561134
rect 379826 525218 380062 525454
rect 380146 525218 380382 525454
rect 379826 524898 380062 525134
rect 380146 524898 380382 525134
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 379826 453218 380062 453454
rect 380146 453218 380382 453454
rect 379826 452898 380062 453134
rect 380146 452898 380382 453134
rect 383546 672938 383782 673174
rect 383866 672938 384102 673174
rect 383546 672618 383782 672854
rect 383866 672618 384102 672854
rect 383546 636938 383782 637174
rect 383866 636938 384102 637174
rect 383546 636618 383782 636854
rect 383866 636618 384102 636854
rect 383546 600938 383782 601174
rect 383866 600938 384102 601174
rect 383546 600618 383782 600854
rect 383866 600618 384102 600854
rect 383546 564938 383782 565174
rect 383866 564938 384102 565174
rect 383546 564618 383782 564854
rect 383866 564618 384102 564854
rect 383546 528938 383782 529174
rect 383866 528938 384102 529174
rect 383546 528618 383782 528854
rect 383866 528618 384102 528854
rect 383546 492938 383782 493174
rect 383866 492938 384102 493174
rect 383546 492618 383782 492854
rect 383866 492618 384102 492854
rect 383546 456938 383782 457174
rect 383866 456938 384102 457174
rect 383546 456618 383782 456854
rect 383866 456618 384102 456854
rect 387266 676658 387502 676894
rect 387586 676658 387822 676894
rect 387266 676338 387502 676574
rect 387586 676338 387822 676574
rect 387266 640658 387502 640894
rect 387586 640658 387822 640894
rect 387266 640338 387502 640574
rect 387586 640338 387822 640574
rect 387266 604658 387502 604894
rect 387586 604658 387822 604894
rect 387266 604338 387502 604574
rect 387586 604338 387822 604574
rect 387266 568658 387502 568894
rect 387586 568658 387822 568894
rect 387266 568338 387502 568574
rect 387586 568338 387822 568574
rect 387266 532658 387502 532894
rect 387586 532658 387822 532894
rect 387266 532338 387502 532574
rect 387586 532338 387822 532574
rect 387266 496658 387502 496894
rect 387586 496658 387822 496894
rect 387266 496338 387502 496574
rect 387586 496338 387822 496574
rect 387266 460658 387502 460894
rect 387586 460658 387822 460894
rect 387266 460338 387502 460574
rect 387586 460338 387822 460574
rect 408986 710362 409222 710598
rect 409306 710362 409542 710598
rect 408986 710042 409222 710278
rect 409306 710042 409542 710278
rect 405266 708442 405502 708678
rect 405586 708442 405822 708678
rect 405266 708122 405502 708358
rect 405586 708122 405822 708358
rect 401546 706522 401782 706758
rect 401866 706522 402102 706758
rect 401546 706202 401782 706438
rect 401866 706202 402102 706438
rect 390986 680378 391222 680614
rect 391306 680378 391542 680614
rect 390986 680058 391222 680294
rect 391306 680058 391542 680294
rect 390986 644378 391222 644614
rect 391306 644378 391542 644614
rect 390986 644058 391222 644294
rect 391306 644058 391542 644294
rect 390986 608378 391222 608614
rect 391306 608378 391542 608614
rect 390986 608058 391222 608294
rect 391306 608058 391542 608294
rect 390986 572378 391222 572614
rect 391306 572378 391542 572614
rect 390986 572058 391222 572294
rect 391306 572058 391542 572294
rect 390986 536378 391222 536614
rect 391306 536378 391542 536614
rect 390986 536058 391222 536294
rect 391306 536058 391542 536294
rect 390986 500378 391222 500614
rect 391306 500378 391542 500614
rect 390986 500058 391222 500294
rect 391306 500058 391542 500294
rect 390986 464378 391222 464614
rect 391306 464378 391542 464614
rect 390986 464058 391222 464294
rect 391306 464058 391542 464294
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 401546 690938 401782 691174
rect 401866 690938 402102 691174
rect 401546 690618 401782 690854
rect 401866 690618 402102 690854
rect 401546 654938 401782 655174
rect 401866 654938 402102 655174
rect 401546 654618 401782 654854
rect 401866 654618 402102 654854
rect 401546 618938 401782 619174
rect 401866 618938 402102 619174
rect 401546 618618 401782 618854
rect 401866 618618 402102 618854
rect 401546 582938 401782 583174
rect 401866 582938 402102 583174
rect 401546 582618 401782 582854
rect 401866 582618 402102 582854
rect 401546 546938 401782 547174
rect 401866 546938 402102 547174
rect 401546 546618 401782 546854
rect 401866 546618 402102 546854
rect 401546 510938 401782 511174
rect 401866 510938 402102 511174
rect 401546 510618 401782 510854
rect 401866 510618 402102 510854
rect 401546 474938 401782 475174
rect 401866 474938 402102 475174
rect 401546 474618 401782 474854
rect 401866 474618 402102 474854
rect 405266 694658 405502 694894
rect 405586 694658 405822 694894
rect 405266 694338 405502 694574
rect 405586 694338 405822 694574
rect 405266 658658 405502 658894
rect 405586 658658 405822 658894
rect 405266 658338 405502 658574
rect 405586 658338 405822 658574
rect 405266 622658 405502 622894
rect 405586 622658 405822 622894
rect 405266 622338 405502 622574
rect 405586 622338 405822 622574
rect 405266 586658 405502 586894
rect 405586 586658 405822 586894
rect 405266 586338 405502 586574
rect 405586 586338 405822 586574
rect 405266 550658 405502 550894
rect 405586 550658 405822 550894
rect 405266 550338 405502 550574
rect 405586 550338 405822 550574
rect 405266 514658 405502 514894
rect 405586 514658 405822 514894
rect 405266 514338 405502 514574
rect 405586 514338 405822 514574
rect 405266 478658 405502 478894
rect 405586 478658 405822 478894
rect 405266 478338 405502 478574
rect 405586 478338 405822 478574
rect 405266 442658 405502 442894
rect 405586 442658 405822 442894
rect 405266 442338 405502 442574
rect 405586 442338 405822 442574
rect 426986 711322 427222 711558
rect 427306 711322 427542 711558
rect 426986 711002 427222 711238
rect 427306 711002 427542 711238
rect 423266 709402 423502 709638
rect 423586 709402 423822 709638
rect 423266 709082 423502 709318
rect 423586 709082 423822 709318
rect 419546 707482 419782 707718
rect 419866 707482 420102 707718
rect 419546 707162 419782 707398
rect 419866 707162 420102 707398
rect 408986 698378 409222 698614
rect 409306 698378 409542 698614
rect 408986 698058 409222 698294
rect 409306 698058 409542 698294
rect 408986 662378 409222 662614
rect 409306 662378 409542 662614
rect 408986 662058 409222 662294
rect 409306 662058 409542 662294
rect 408986 626378 409222 626614
rect 409306 626378 409542 626614
rect 408986 626058 409222 626294
rect 409306 626058 409542 626294
rect 408986 590378 409222 590614
rect 409306 590378 409542 590614
rect 408986 590058 409222 590294
rect 409306 590058 409542 590294
rect 408986 554378 409222 554614
rect 409306 554378 409542 554614
rect 408986 554058 409222 554294
rect 409306 554058 409542 554294
rect 408986 518378 409222 518614
rect 409306 518378 409542 518614
rect 408986 518058 409222 518294
rect 409306 518058 409542 518294
rect 408986 482378 409222 482614
rect 409306 482378 409542 482614
rect 408986 482058 409222 482294
rect 409306 482058 409542 482294
rect 408986 446378 409222 446614
rect 409306 446378 409542 446614
rect 408986 446058 409222 446294
rect 409306 446058 409542 446294
rect 415826 705562 416062 705798
rect 416146 705562 416382 705798
rect 415826 705242 416062 705478
rect 416146 705242 416382 705478
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 415826 561218 416062 561454
rect 416146 561218 416382 561454
rect 415826 560898 416062 561134
rect 416146 560898 416382 561134
rect 415826 525218 416062 525454
rect 416146 525218 416382 525454
rect 415826 524898 416062 525134
rect 416146 524898 416382 525134
rect 415826 489218 416062 489454
rect 416146 489218 416382 489454
rect 415826 488898 416062 489134
rect 416146 488898 416382 489134
rect 415826 453218 416062 453454
rect 416146 453218 416382 453454
rect 415826 452898 416062 453134
rect 416146 452898 416382 453134
rect 419546 672938 419782 673174
rect 419866 672938 420102 673174
rect 419546 672618 419782 672854
rect 419866 672618 420102 672854
rect 419546 636938 419782 637174
rect 419866 636938 420102 637174
rect 419546 636618 419782 636854
rect 419866 636618 420102 636854
rect 419546 600938 419782 601174
rect 419866 600938 420102 601174
rect 419546 600618 419782 600854
rect 419866 600618 420102 600854
rect 419546 564938 419782 565174
rect 419866 564938 420102 565174
rect 419546 564618 419782 564854
rect 419866 564618 420102 564854
rect 419546 528938 419782 529174
rect 419866 528938 420102 529174
rect 419546 528618 419782 528854
rect 419866 528618 420102 528854
rect 419546 492938 419782 493174
rect 419866 492938 420102 493174
rect 419546 492618 419782 492854
rect 419866 492618 420102 492854
rect 419546 456938 419782 457174
rect 419866 456938 420102 457174
rect 419546 456618 419782 456854
rect 419866 456618 420102 456854
rect 423266 676658 423502 676894
rect 423586 676658 423822 676894
rect 423266 676338 423502 676574
rect 423586 676338 423822 676574
rect 423266 640658 423502 640894
rect 423586 640658 423822 640894
rect 423266 640338 423502 640574
rect 423586 640338 423822 640574
rect 423266 604658 423502 604894
rect 423586 604658 423822 604894
rect 423266 604338 423502 604574
rect 423586 604338 423822 604574
rect 423266 568658 423502 568894
rect 423586 568658 423822 568894
rect 423266 568338 423502 568574
rect 423586 568338 423822 568574
rect 423266 532658 423502 532894
rect 423586 532658 423822 532894
rect 423266 532338 423502 532574
rect 423586 532338 423822 532574
rect 423266 496658 423502 496894
rect 423586 496658 423822 496894
rect 423266 496338 423502 496574
rect 423586 496338 423822 496574
rect 423266 460658 423502 460894
rect 423586 460658 423822 460894
rect 423266 460338 423502 460574
rect 423586 460338 423822 460574
rect 444986 710362 445222 710598
rect 445306 710362 445542 710598
rect 444986 710042 445222 710278
rect 445306 710042 445542 710278
rect 441266 708442 441502 708678
rect 441586 708442 441822 708678
rect 441266 708122 441502 708358
rect 441586 708122 441822 708358
rect 437546 706522 437782 706758
rect 437866 706522 438102 706758
rect 437546 706202 437782 706438
rect 437866 706202 438102 706438
rect 426986 680378 427222 680614
rect 427306 680378 427542 680614
rect 426986 680058 427222 680294
rect 427306 680058 427542 680294
rect 426986 644378 427222 644614
rect 427306 644378 427542 644614
rect 426986 644058 427222 644294
rect 427306 644058 427542 644294
rect 426986 608378 427222 608614
rect 427306 608378 427542 608614
rect 426986 608058 427222 608294
rect 427306 608058 427542 608294
rect 426986 572378 427222 572614
rect 427306 572378 427542 572614
rect 426986 572058 427222 572294
rect 427306 572058 427542 572294
rect 426986 536378 427222 536614
rect 427306 536378 427542 536614
rect 426986 536058 427222 536294
rect 427306 536058 427542 536294
rect 426986 500378 427222 500614
rect 427306 500378 427542 500614
rect 426986 500058 427222 500294
rect 427306 500058 427542 500294
rect 426986 464378 427222 464614
rect 427306 464378 427542 464614
rect 426986 464058 427222 464294
rect 427306 464058 427542 464294
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 437546 690938 437782 691174
rect 437866 690938 438102 691174
rect 437546 690618 437782 690854
rect 437866 690618 438102 690854
rect 437546 654938 437782 655174
rect 437866 654938 438102 655174
rect 437546 654618 437782 654854
rect 437866 654618 438102 654854
rect 437546 618938 437782 619174
rect 437866 618938 438102 619174
rect 437546 618618 437782 618854
rect 437866 618618 438102 618854
rect 437546 582938 437782 583174
rect 437866 582938 438102 583174
rect 437546 582618 437782 582854
rect 437866 582618 438102 582854
rect 437546 546938 437782 547174
rect 437866 546938 438102 547174
rect 437546 546618 437782 546854
rect 437866 546618 438102 546854
rect 437546 510938 437782 511174
rect 437866 510938 438102 511174
rect 437546 510618 437782 510854
rect 437866 510618 438102 510854
rect 437546 474938 437782 475174
rect 437866 474938 438102 475174
rect 437546 474618 437782 474854
rect 437866 474618 438102 474854
rect 441266 694658 441502 694894
rect 441586 694658 441822 694894
rect 441266 694338 441502 694574
rect 441586 694338 441822 694574
rect 441266 658658 441502 658894
rect 441586 658658 441822 658894
rect 441266 658338 441502 658574
rect 441586 658338 441822 658574
rect 441266 622658 441502 622894
rect 441586 622658 441822 622894
rect 441266 622338 441502 622574
rect 441586 622338 441822 622574
rect 441266 586658 441502 586894
rect 441586 586658 441822 586894
rect 441266 586338 441502 586574
rect 441586 586338 441822 586574
rect 441266 550658 441502 550894
rect 441586 550658 441822 550894
rect 441266 550338 441502 550574
rect 441586 550338 441822 550574
rect 441266 514658 441502 514894
rect 441586 514658 441822 514894
rect 441266 514338 441502 514574
rect 441586 514338 441822 514574
rect 441266 478658 441502 478894
rect 441586 478658 441822 478894
rect 441266 478338 441502 478574
rect 441586 478338 441822 478574
rect 441266 442658 441502 442894
rect 441586 442658 441822 442894
rect 441266 442338 441502 442574
rect 441586 442338 441822 442574
rect 462986 711322 463222 711558
rect 463306 711322 463542 711558
rect 462986 711002 463222 711238
rect 463306 711002 463542 711238
rect 459266 709402 459502 709638
rect 459586 709402 459822 709638
rect 459266 709082 459502 709318
rect 459586 709082 459822 709318
rect 455546 707482 455782 707718
rect 455866 707482 456102 707718
rect 455546 707162 455782 707398
rect 455866 707162 456102 707398
rect 444986 698378 445222 698614
rect 445306 698378 445542 698614
rect 444986 698058 445222 698294
rect 445306 698058 445542 698294
rect 444986 662378 445222 662614
rect 445306 662378 445542 662614
rect 444986 662058 445222 662294
rect 445306 662058 445542 662294
rect 444986 626378 445222 626614
rect 445306 626378 445542 626614
rect 444986 626058 445222 626294
rect 445306 626058 445542 626294
rect 444986 590378 445222 590614
rect 445306 590378 445542 590614
rect 444986 590058 445222 590294
rect 445306 590058 445542 590294
rect 444986 554378 445222 554614
rect 445306 554378 445542 554614
rect 444986 554058 445222 554294
rect 445306 554058 445542 554294
rect 444986 518378 445222 518614
rect 445306 518378 445542 518614
rect 444986 518058 445222 518294
rect 445306 518058 445542 518294
rect 444986 482378 445222 482614
rect 445306 482378 445542 482614
rect 444986 482058 445222 482294
rect 445306 482058 445542 482294
rect 444986 446378 445222 446614
rect 445306 446378 445542 446614
rect 444986 446058 445222 446294
rect 445306 446058 445542 446294
rect 451826 705562 452062 705798
rect 452146 705562 452382 705798
rect 451826 705242 452062 705478
rect 452146 705242 452382 705478
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 451826 453218 452062 453454
rect 452146 453218 452382 453454
rect 451826 452898 452062 453134
rect 452146 452898 452382 453134
rect 455546 672938 455782 673174
rect 455866 672938 456102 673174
rect 455546 672618 455782 672854
rect 455866 672618 456102 672854
rect 455546 636938 455782 637174
rect 455866 636938 456102 637174
rect 455546 636618 455782 636854
rect 455866 636618 456102 636854
rect 455546 600938 455782 601174
rect 455866 600938 456102 601174
rect 455546 600618 455782 600854
rect 455866 600618 456102 600854
rect 455546 564938 455782 565174
rect 455866 564938 456102 565174
rect 455546 564618 455782 564854
rect 455866 564618 456102 564854
rect 455546 528938 455782 529174
rect 455866 528938 456102 529174
rect 455546 528618 455782 528854
rect 455866 528618 456102 528854
rect 455546 492938 455782 493174
rect 455866 492938 456102 493174
rect 455546 492618 455782 492854
rect 455866 492618 456102 492854
rect 455546 456938 455782 457174
rect 455866 456938 456102 457174
rect 455546 456618 455782 456854
rect 455866 456618 456102 456854
rect 459266 676658 459502 676894
rect 459586 676658 459822 676894
rect 459266 676338 459502 676574
rect 459586 676338 459822 676574
rect 459266 640658 459502 640894
rect 459586 640658 459822 640894
rect 459266 640338 459502 640574
rect 459586 640338 459822 640574
rect 459266 604658 459502 604894
rect 459586 604658 459822 604894
rect 459266 604338 459502 604574
rect 459586 604338 459822 604574
rect 459266 568658 459502 568894
rect 459586 568658 459822 568894
rect 459266 568338 459502 568574
rect 459586 568338 459822 568574
rect 459266 532658 459502 532894
rect 459586 532658 459822 532894
rect 459266 532338 459502 532574
rect 459586 532338 459822 532574
rect 459266 496658 459502 496894
rect 459586 496658 459822 496894
rect 459266 496338 459502 496574
rect 459586 496338 459822 496574
rect 459266 460658 459502 460894
rect 459586 460658 459822 460894
rect 459266 460338 459502 460574
rect 459586 460338 459822 460574
rect 480986 710362 481222 710598
rect 481306 710362 481542 710598
rect 480986 710042 481222 710278
rect 481306 710042 481542 710278
rect 477266 708442 477502 708678
rect 477586 708442 477822 708678
rect 477266 708122 477502 708358
rect 477586 708122 477822 708358
rect 473546 706522 473782 706758
rect 473866 706522 474102 706758
rect 473546 706202 473782 706438
rect 473866 706202 474102 706438
rect 462986 680378 463222 680614
rect 463306 680378 463542 680614
rect 462986 680058 463222 680294
rect 463306 680058 463542 680294
rect 462986 644378 463222 644614
rect 463306 644378 463542 644614
rect 462986 644058 463222 644294
rect 463306 644058 463542 644294
rect 462986 608378 463222 608614
rect 463306 608378 463542 608614
rect 462986 608058 463222 608294
rect 463306 608058 463542 608294
rect 462986 572378 463222 572614
rect 463306 572378 463542 572614
rect 462986 572058 463222 572294
rect 463306 572058 463542 572294
rect 462986 536378 463222 536614
rect 463306 536378 463542 536614
rect 462986 536058 463222 536294
rect 463306 536058 463542 536294
rect 462986 500378 463222 500614
rect 463306 500378 463542 500614
rect 462986 500058 463222 500294
rect 463306 500058 463542 500294
rect 462986 464378 463222 464614
rect 463306 464378 463542 464614
rect 462986 464058 463222 464294
rect 463306 464058 463542 464294
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 473546 690938 473782 691174
rect 473866 690938 474102 691174
rect 473546 690618 473782 690854
rect 473866 690618 474102 690854
rect 473546 654938 473782 655174
rect 473866 654938 474102 655174
rect 473546 654618 473782 654854
rect 473866 654618 474102 654854
rect 473546 618938 473782 619174
rect 473866 618938 474102 619174
rect 473546 618618 473782 618854
rect 473866 618618 474102 618854
rect 473546 582938 473782 583174
rect 473866 582938 474102 583174
rect 473546 582618 473782 582854
rect 473866 582618 474102 582854
rect 473546 546938 473782 547174
rect 473866 546938 474102 547174
rect 473546 546618 473782 546854
rect 473866 546618 474102 546854
rect 473546 510938 473782 511174
rect 473866 510938 474102 511174
rect 473546 510618 473782 510854
rect 473866 510618 474102 510854
rect 473546 474938 473782 475174
rect 473866 474938 474102 475174
rect 473546 474618 473782 474854
rect 473866 474618 474102 474854
rect 477266 694658 477502 694894
rect 477586 694658 477822 694894
rect 477266 694338 477502 694574
rect 477586 694338 477822 694574
rect 477266 658658 477502 658894
rect 477586 658658 477822 658894
rect 477266 658338 477502 658574
rect 477586 658338 477822 658574
rect 477266 622658 477502 622894
rect 477586 622658 477822 622894
rect 477266 622338 477502 622574
rect 477586 622338 477822 622574
rect 477266 586658 477502 586894
rect 477586 586658 477822 586894
rect 477266 586338 477502 586574
rect 477586 586338 477822 586574
rect 477266 550658 477502 550894
rect 477586 550658 477822 550894
rect 477266 550338 477502 550574
rect 477586 550338 477822 550574
rect 477266 514658 477502 514894
rect 477586 514658 477822 514894
rect 477266 514338 477502 514574
rect 477586 514338 477822 514574
rect 477266 478658 477502 478894
rect 477586 478658 477822 478894
rect 477266 478338 477502 478574
rect 477586 478338 477822 478574
rect 477266 442658 477502 442894
rect 477586 442658 477822 442894
rect 477266 442338 477502 442574
rect 477586 442338 477822 442574
rect 498986 711322 499222 711558
rect 499306 711322 499542 711558
rect 498986 711002 499222 711238
rect 499306 711002 499542 711238
rect 495266 709402 495502 709638
rect 495586 709402 495822 709638
rect 495266 709082 495502 709318
rect 495586 709082 495822 709318
rect 491546 707482 491782 707718
rect 491866 707482 492102 707718
rect 491546 707162 491782 707398
rect 491866 707162 492102 707398
rect 480986 698378 481222 698614
rect 481306 698378 481542 698614
rect 480986 698058 481222 698294
rect 481306 698058 481542 698294
rect 480986 662378 481222 662614
rect 481306 662378 481542 662614
rect 480986 662058 481222 662294
rect 481306 662058 481542 662294
rect 480986 626378 481222 626614
rect 481306 626378 481542 626614
rect 480986 626058 481222 626294
rect 481306 626058 481542 626294
rect 480986 590378 481222 590614
rect 481306 590378 481542 590614
rect 480986 590058 481222 590294
rect 481306 590058 481542 590294
rect 480986 554378 481222 554614
rect 481306 554378 481542 554614
rect 480986 554058 481222 554294
rect 481306 554058 481542 554294
rect 480986 518378 481222 518614
rect 481306 518378 481542 518614
rect 480986 518058 481222 518294
rect 481306 518058 481542 518294
rect 480986 482378 481222 482614
rect 481306 482378 481542 482614
rect 480986 482058 481222 482294
rect 481306 482058 481542 482294
rect 480986 446378 481222 446614
rect 481306 446378 481542 446614
rect 480986 446058 481222 446294
rect 481306 446058 481542 446294
rect 487826 705562 488062 705798
rect 488146 705562 488382 705798
rect 487826 705242 488062 705478
rect 488146 705242 488382 705478
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 487826 453218 488062 453454
rect 488146 453218 488382 453454
rect 487826 452898 488062 453134
rect 488146 452898 488382 453134
rect 244250 435218 244486 435454
rect 244250 434898 244486 435134
rect 274970 435218 275206 435454
rect 274970 434898 275206 435134
rect 305690 435218 305926 435454
rect 305690 434898 305926 435134
rect 336410 435218 336646 435454
rect 336410 434898 336646 435134
rect 367130 435218 367366 435454
rect 367130 434898 367366 435134
rect 397850 435218 398086 435454
rect 397850 434898 398086 435134
rect 428570 435218 428806 435454
rect 428570 434898 428806 435134
rect 459290 435218 459526 435454
rect 459290 434898 459526 435134
rect 490010 435218 490246 435454
rect 490010 434898 490246 435134
rect 259610 417218 259846 417454
rect 259610 416898 259846 417134
rect 290330 417218 290566 417454
rect 290330 416898 290566 417134
rect 321050 417218 321286 417454
rect 321050 416898 321286 417134
rect 351770 417218 352006 417454
rect 351770 416898 352006 417134
rect 382490 417218 382726 417454
rect 382490 416898 382726 417134
rect 413210 417218 413446 417454
rect 413210 416898 413446 417134
rect 443930 417218 444166 417454
rect 443930 416898 444166 417134
rect 474650 417218 474886 417454
rect 474650 416898 474886 417134
rect 244250 399218 244486 399454
rect 244250 398898 244486 399134
rect 274970 399218 275206 399454
rect 274970 398898 275206 399134
rect 305690 399218 305926 399454
rect 305690 398898 305926 399134
rect 336410 399218 336646 399454
rect 336410 398898 336646 399134
rect 367130 399218 367366 399454
rect 367130 398898 367366 399134
rect 397850 399218 398086 399454
rect 397850 398898 398086 399134
rect 428570 399218 428806 399454
rect 428570 398898 428806 399134
rect 459290 399218 459526 399454
rect 459290 398898 459526 399134
rect 490010 399218 490246 399454
rect 490010 398898 490246 399134
rect 259610 381218 259846 381454
rect 259610 380898 259846 381134
rect 290330 381218 290566 381454
rect 290330 380898 290566 381134
rect 321050 381218 321286 381454
rect 321050 380898 321286 381134
rect 351770 381218 352006 381454
rect 351770 380898 352006 381134
rect 382490 381218 382726 381454
rect 382490 380898 382726 381134
rect 413210 381218 413446 381454
rect 413210 380898 413446 381134
rect 443930 381218 444166 381454
rect 443930 380898 444166 381134
rect 474650 381218 474886 381454
rect 474650 380898 474886 381134
rect 244250 363218 244486 363454
rect 244250 362898 244486 363134
rect 274970 363218 275206 363454
rect 274970 362898 275206 363134
rect 305690 363218 305926 363454
rect 305690 362898 305926 363134
rect 336410 363218 336646 363454
rect 336410 362898 336646 363134
rect 367130 363218 367366 363454
rect 367130 362898 367366 363134
rect 397850 363218 398086 363454
rect 397850 362898 398086 363134
rect 428570 363218 428806 363454
rect 428570 362898 428806 363134
rect 459290 363218 459526 363454
rect 459290 362898 459526 363134
rect 490010 363218 490246 363454
rect 490010 362898 490246 363134
rect 259610 345218 259846 345454
rect 259610 344898 259846 345134
rect 290330 345218 290566 345454
rect 290330 344898 290566 345134
rect 321050 345218 321286 345454
rect 321050 344898 321286 345134
rect 351770 345218 352006 345454
rect 351770 344898 352006 345134
rect 382490 345218 382726 345454
rect 382490 344898 382726 345134
rect 413210 345218 413446 345454
rect 413210 344898 413446 345134
rect 443930 345218 444166 345454
rect 443930 344898 444166 345134
rect 474650 345218 474886 345454
rect 474650 344898 474886 345134
rect 244250 327218 244486 327454
rect 244250 326898 244486 327134
rect 274970 327218 275206 327454
rect 274970 326898 275206 327134
rect 305690 327218 305926 327454
rect 305690 326898 305926 327134
rect 336410 327218 336646 327454
rect 336410 326898 336646 327134
rect 367130 327218 367366 327454
rect 367130 326898 367366 327134
rect 397850 327218 398086 327454
rect 397850 326898 398086 327134
rect 428570 327218 428806 327454
rect 428570 326898 428806 327134
rect 459290 327218 459526 327454
rect 459290 326898 459526 327134
rect 490010 327218 490246 327454
rect 490010 326898 490246 327134
rect 259610 309218 259846 309454
rect 259610 308898 259846 309134
rect 290330 309218 290566 309454
rect 290330 308898 290566 309134
rect 321050 309218 321286 309454
rect 321050 308898 321286 309134
rect 351770 309218 352006 309454
rect 351770 308898 352006 309134
rect 382490 309218 382726 309454
rect 382490 308898 382726 309134
rect 413210 309218 413446 309454
rect 413210 308898 413446 309134
rect 443930 309218 444166 309454
rect 443930 308898 444166 309134
rect 474650 309218 474886 309454
rect 474650 308898 474886 309134
rect 244250 291218 244486 291454
rect 244250 290898 244486 291134
rect 274970 291218 275206 291454
rect 274970 290898 275206 291134
rect 305690 291218 305926 291454
rect 305690 290898 305926 291134
rect 336410 291218 336646 291454
rect 336410 290898 336646 291134
rect 367130 291218 367366 291454
rect 367130 290898 367366 291134
rect 397850 291218 398086 291454
rect 397850 290898 398086 291134
rect 428570 291218 428806 291454
rect 428570 290898 428806 291134
rect 459290 291218 459526 291454
rect 459290 290898 459526 291134
rect 490010 291218 490246 291454
rect 490010 290898 490246 291134
rect 259610 273218 259846 273454
rect 259610 272898 259846 273134
rect 290330 273218 290566 273454
rect 290330 272898 290566 273134
rect 321050 273218 321286 273454
rect 321050 272898 321286 273134
rect 351770 273218 352006 273454
rect 351770 272898 352006 273134
rect 382490 273218 382726 273454
rect 382490 272898 382726 273134
rect 413210 273218 413446 273454
rect 413210 272898 413446 273134
rect 443930 273218 444166 273454
rect 443930 272898 444166 273134
rect 474650 273218 474886 273454
rect 474650 272898 474886 273134
rect 244250 255218 244486 255454
rect 244250 254898 244486 255134
rect 274970 255218 275206 255454
rect 274970 254898 275206 255134
rect 305690 255218 305926 255454
rect 305690 254898 305926 255134
rect 336410 255218 336646 255454
rect 336410 254898 336646 255134
rect 367130 255218 367366 255454
rect 367130 254898 367366 255134
rect 397850 255218 398086 255454
rect 397850 254898 398086 255134
rect 428570 255218 428806 255454
rect 428570 254898 428806 255134
rect 459290 255218 459526 255454
rect 459290 254898 459526 255134
rect 490010 255218 490246 255454
rect 490010 254898 490246 255134
rect 259610 237218 259846 237454
rect 259610 236898 259846 237134
rect 290330 237218 290566 237454
rect 290330 236898 290566 237134
rect 321050 237218 321286 237454
rect 321050 236898 321286 237134
rect 351770 237218 352006 237454
rect 351770 236898 352006 237134
rect 382490 237218 382726 237454
rect 382490 236898 382726 237134
rect 413210 237218 413446 237454
rect 413210 236898 413446 237134
rect 443930 237218 444166 237454
rect 443930 236898 444166 237134
rect 474650 237218 474886 237454
rect 474650 236898 474886 237134
rect 244250 219218 244486 219454
rect 244250 218898 244486 219134
rect 274970 219218 275206 219454
rect 274970 218898 275206 219134
rect 305690 219218 305926 219454
rect 305690 218898 305926 219134
rect 336410 219218 336646 219454
rect 336410 218898 336646 219134
rect 367130 219218 367366 219454
rect 367130 218898 367366 219134
rect 397850 219218 398086 219454
rect 397850 218898 398086 219134
rect 428570 219218 428806 219454
rect 428570 218898 428806 219134
rect 459290 219218 459526 219454
rect 459290 218898 459526 219134
rect 490010 219218 490246 219454
rect 490010 218898 490246 219134
rect 259610 201218 259846 201454
rect 259610 200898 259846 201134
rect 290330 201218 290566 201454
rect 290330 200898 290566 201134
rect 321050 201218 321286 201454
rect 321050 200898 321286 201134
rect 351770 201218 352006 201454
rect 351770 200898 352006 201134
rect 382490 201218 382726 201454
rect 382490 200898 382726 201134
rect 413210 201218 413446 201454
rect 413210 200898 413446 201134
rect 443930 201218 444166 201454
rect 443930 200898 444166 201134
rect 474650 201218 474886 201454
rect 474650 200898 474886 201134
rect 244250 183218 244486 183454
rect 244250 182898 244486 183134
rect 274970 183218 275206 183454
rect 274970 182898 275206 183134
rect 305690 183218 305926 183454
rect 305690 182898 305926 183134
rect 336410 183218 336646 183454
rect 336410 182898 336646 183134
rect 367130 183218 367366 183454
rect 367130 182898 367366 183134
rect 397850 183218 398086 183454
rect 397850 182898 398086 183134
rect 428570 183218 428806 183454
rect 428570 182898 428806 183134
rect 459290 183218 459526 183454
rect 459290 182898 459526 183134
rect 490010 183218 490246 183454
rect 490010 182898 490246 183134
rect 491546 672938 491782 673174
rect 491866 672938 492102 673174
rect 491546 672618 491782 672854
rect 491866 672618 492102 672854
rect 491546 636938 491782 637174
rect 491866 636938 492102 637174
rect 491546 636618 491782 636854
rect 491866 636618 492102 636854
rect 491546 600938 491782 601174
rect 491866 600938 492102 601174
rect 491546 600618 491782 600854
rect 491866 600618 492102 600854
rect 491546 564938 491782 565174
rect 491866 564938 492102 565174
rect 491546 564618 491782 564854
rect 491866 564618 492102 564854
rect 491546 528938 491782 529174
rect 491866 528938 492102 529174
rect 491546 528618 491782 528854
rect 491866 528618 492102 528854
rect 491546 492938 491782 493174
rect 491866 492938 492102 493174
rect 491546 492618 491782 492854
rect 491866 492618 492102 492854
rect 491546 456938 491782 457174
rect 491866 456938 492102 457174
rect 491546 456618 491782 456854
rect 491866 456618 492102 456854
rect 495266 676658 495502 676894
rect 495586 676658 495822 676894
rect 495266 676338 495502 676574
rect 495586 676338 495822 676574
rect 495266 640658 495502 640894
rect 495586 640658 495822 640894
rect 495266 640338 495502 640574
rect 495586 640338 495822 640574
rect 495266 604658 495502 604894
rect 495586 604658 495822 604894
rect 495266 604338 495502 604574
rect 495586 604338 495822 604574
rect 495266 568658 495502 568894
rect 495586 568658 495822 568894
rect 495266 568338 495502 568574
rect 495586 568338 495822 568574
rect 495266 532658 495502 532894
rect 495586 532658 495822 532894
rect 495266 532338 495502 532574
rect 495586 532338 495822 532574
rect 495266 496658 495502 496894
rect 495586 496658 495822 496894
rect 495266 496338 495502 496574
rect 495586 496338 495822 496574
rect 495266 460658 495502 460894
rect 495586 460658 495822 460894
rect 495266 460338 495502 460574
rect 495586 460338 495822 460574
rect 516986 710362 517222 710598
rect 517306 710362 517542 710598
rect 516986 710042 517222 710278
rect 517306 710042 517542 710278
rect 513266 708442 513502 708678
rect 513586 708442 513822 708678
rect 513266 708122 513502 708358
rect 513586 708122 513822 708358
rect 509546 706522 509782 706758
rect 509866 706522 510102 706758
rect 509546 706202 509782 706438
rect 509866 706202 510102 706438
rect 498986 680378 499222 680614
rect 499306 680378 499542 680614
rect 498986 680058 499222 680294
rect 499306 680058 499542 680294
rect 498986 644378 499222 644614
rect 499306 644378 499542 644614
rect 498986 644058 499222 644294
rect 499306 644058 499542 644294
rect 498986 608378 499222 608614
rect 499306 608378 499542 608614
rect 498986 608058 499222 608294
rect 499306 608058 499542 608294
rect 498986 572378 499222 572614
rect 499306 572378 499542 572614
rect 498986 572058 499222 572294
rect 499306 572058 499542 572294
rect 498986 536378 499222 536614
rect 499306 536378 499542 536614
rect 498986 536058 499222 536294
rect 499306 536058 499542 536294
rect 498986 500378 499222 500614
rect 499306 500378 499542 500614
rect 498986 500058 499222 500294
rect 499306 500058 499542 500294
rect 498986 464378 499222 464614
rect 499306 464378 499542 464614
rect 498986 464058 499222 464294
rect 499306 464058 499542 464294
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 235826 165218 236062 165454
rect 236146 165218 236382 165454
rect 235826 164898 236062 165134
rect 236146 164898 236382 165134
rect 235826 129218 236062 129454
rect 236146 129218 236382 129454
rect 235826 128898 236062 129134
rect 236146 128898 236382 129134
rect 235826 93218 236062 93454
rect 236146 93218 236382 93454
rect 235826 92898 236062 93134
rect 236146 92898 236382 93134
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -1542 236062 -1306
rect 236146 -1542 236382 -1306
rect 235826 -1862 236062 -1626
rect 236146 -1862 236382 -1626
rect 239546 168938 239782 169174
rect 239866 168938 240102 169174
rect 239546 168618 239782 168854
rect 239866 168618 240102 168854
rect 239546 132938 239782 133174
rect 239866 132938 240102 133174
rect 239546 132618 239782 132854
rect 239866 132618 240102 132854
rect 239546 96938 239782 97174
rect 239866 96938 240102 97174
rect 239546 96618 239782 96854
rect 239866 96618 240102 96854
rect 239546 60938 239782 61174
rect 239866 60938 240102 61174
rect 239546 60618 239782 60854
rect 239866 60618 240102 60854
rect 239546 24938 239782 25174
rect 239866 24938 240102 25174
rect 239546 24618 239782 24854
rect 239866 24618 240102 24854
rect 239546 -3462 239782 -3226
rect 239866 -3462 240102 -3226
rect 239546 -3782 239782 -3546
rect 239866 -3782 240102 -3546
rect 243266 172658 243502 172894
rect 243586 172658 243822 172894
rect 243266 172338 243502 172574
rect 243586 172338 243822 172574
rect 243266 136658 243502 136894
rect 243586 136658 243822 136894
rect 243266 136338 243502 136574
rect 243586 136338 243822 136574
rect 243266 100658 243502 100894
rect 243586 100658 243822 100894
rect 243266 100338 243502 100574
rect 243586 100338 243822 100574
rect 243266 64658 243502 64894
rect 243586 64658 243822 64894
rect 243266 64338 243502 64574
rect 243586 64338 243822 64574
rect 243266 28658 243502 28894
rect 243586 28658 243822 28894
rect 243266 28338 243502 28574
rect 243586 28338 243822 28574
rect 243266 -5382 243502 -5146
rect 243586 -5382 243822 -5146
rect 243266 -5702 243502 -5466
rect 243586 -5702 243822 -5466
rect 246986 176378 247222 176614
rect 247306 176378 247542 176614
rect 246986 176058 247222 176294
rect 247306 176058 247542 176294
rect 246986 140378 247222 140614
rect 247306 140378 247542 140614
rect 246986 140058 247222 140294
rect 247306 140058 247542 140294
rect 246986 104378 247222 104614
rect 247306 104378 247542 104614
rect 246986 104058 247222 104294
rect 247306 104058 247542 104294
rect 246986 68378 247222 68614
rect 247306 68378 247542 68614
rect 246986 68058 247222 68294
rect 247306 68058 247542 68294
rect 246986 32378 247222 32614
rect 247306 32378 247542 32614
rect 246986 32058 247222 32294
rect 247306 32058 247542 32294
rect 228986 -6342 229222 -6106
rect 229306 -6342 229542 -6106
rect 228986 -6662 229222 -6426
rect 229306 -6662 229542 -6426
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 253826 111218 254062 111454
rect 254146 111218 254382 111454
rect 253826 110898 254062 111134
rect 254146 110898 254382 111134
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 257546 150938 257782 151174
rect 257866 150938 258102 151174
rect 257546 150618 257782 150854
rect 257866 150618 258102 150854
rect 257546 114938 257782 115174
rect 257866 114938 258102 115174
rect 257546 114618 257782 114854
rect 257866 114618 258102 114854
rect 257546 78938 257782 79174
rect 257866 78938 258102 79174
rect 257546 78618 257782 78854
rect 257866 78618 258102 78854
rect 257546 42938 257782 43174
rect 257866 42938 258102 43174
rect 257546 42618 257782 42854
rect 257866 42618 258102 42854
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 257546 -2502 257782 -2266
rect 257866 -2502 258102 -2266
rect 257546 -2822 257782 -2586
rect 257866 -2822 258102 -2586
rect 261266 154658 261502 154894
rect 261586 154658 261822 154894
rect 261266 154338 261502 154574
rect 261586 154338 261822 154574
rect 261266 118658 261502 118894
rect 261586 118658 261822 118894
rect 261266 118338 261502 118574
rect 261586 118338 261822 118574
rect 261266 82658 261502 82894
rect 261586 82658 261822 82894
rect 261266 82338 261502 82574
rect 261586 82338 261822 82574
rect 261266 46658 261502 46894
rect 261586 46658 261822 46894
rect 261266 46338 261502 46574
rect 261586 46338 261822 46574
rect 261266 10658 261502 10894
rect 261586 10658 261822 10894
rect 261266 10338 261502 10574
rect 261586 10338 261822 10574
rect 261266 -4422 261502 -4186
rect 261586 -4422 261822 -4186
rect 261266 -4742 261502 -4506
rect 261586 -4742 261822 -4506
rect 264986 158378 265222 158614
rect 265306 158378 265542 158614
rect 264986 158058 265222 158294
rect 265306 158058 265542 158294
rect 264986 122378 265222 122614
rect 265306 122378 265542 122614
rect 264986 122058 265222 122294
rect 265306 122058 265542 122294
rect 264986 86378 265222 86614
rect 265306 86378 265542 86614
rect 264986 86058 265222 86294
rect 265306 86058 265542 86294
rect 264986 50378 265222 50614
rect 265306 50378 265542 50614
rect 264986 50058 265222 50294
rect 265306 50058 265542 50294
rect 264986 14378 265222 14614
rect 265306 14378 265542 14614
rect 264986 14058 265222 14294
rect 265306 14058 265542 14294
rect 246986 -7302 247222 -7066
rect 247306 -7302 247542 -7066
rect 246986 -7622 247222 -7386
rect 247306 -7622 247542 -7386
rect 271826 165218 272062 165454
rect 272146 165218 272382 165454
rect 271826 164898 272062 165134
rect 272146 164898 272382 165134
rect 271826 129218 272062 129454
rect 272146 129218 272382 129454
rect 271826 128898 272062 129134
rect 272146 128898 272382 129134
rect 271826 93218 272062 93454
rect 272146 93218 272382 93454
rect 271826 92898 272062 93134
rect 272146 92898 272382 93134
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -1542 272062 -1306
rect 272146 -1542 272382 -1306
rect 271826 -1862 272062 -1626
rect 272146 -1862 272382 -1626
rect 275546 168938 275782 169174
rect 275866 168938 276102 169174
rect 275546 168618 275782 168854
rect 275866 168618 276102 168854
rect 275546 132938 275782 133174
rect 275866 132938 276102 133174
rect 275546 132618 275782 132854
rect 275866 132618 276102 132854
rect 275546 96938 275782 97174
rect 275866 96938 276102 97174
rect 275546 96618 275782 96854
rect 275866 96618 276102 96854
rect 275546 60938 275782 61174
rect 275866 60938 276102 61174
rect 275546 60618 275782 60854
rect 275866 60618 276102 60854
rect 275546 24938 275782 25174
rect 275866 24938 276102 25174
rect 275546 24618 275782 24854
rect 275866 24618 276102 24854
rect 275546 -3462 275782 -3226
rect 275866 -3462 276102 -3226
rect 275546 -3782 275782 -3546
rect 275866 -3782 276102 -3546
rect 279266 172658 279502 172894
rect 279586 172658 279822 172894
rect 279266 172338 279502 172574
rect 279586 172338 279822 172574
rect 279266 136658 279502 136894
rect 279586 136658 279822 136894
rect 279266 136338 279502 136574
rect 279586 136338 279822 136574
rect 279266 100658 279502 100894
rect 279586 100658 279822 100894
rect 279266 100338 279502 100574
rect 279586 100338 279822 100574
rect 279266 64658 279502 64894
rect 279586 64658 279822 64894
rect 279266 64338 279502 64574
rect 279586 64338 279822 64574
rect 279266 28658 279502 28894
rect 279586 28658 279822 28894
rect 279266 28338 279502 28574
rect 279586 28338 279822 28574
rect 279266 -5382 279502 -5146
rect 279586 -5382 279822 -5146
rect 279266 -5702 279502 -5466
rect 279586 -5702 279822 -5466
rect 282986 176378 283222 176614
rect 283306 176378 283542 176614
rect 282986 176058 283222 176294
rect 283306 176058 283542 176294
rect 282986 140378 283222 140614
rect 283306 140378 283542 140614
rect 282986 140058 283222 140294
rect 283306 140058 283542 140294
rect 282986 104378 283222 104614
rect 283306 104378 283542 104614
rect 282986 104058 283222 104294
rect 283306 104058 283542 104294
rect 282986 68378 283222 68614
rect 283306 68378 283542 68614
rect 282986 68058 283222 68294
rect 283306 68058 283542 68294
rect 282986 32378 283222 32614
rect 283306 32378 283542 32614
rect 282986 32058 283222 32294
rect 283306 32058 283542 32294
rect 264986 -6342 265222 -6106
rect 265306 -6342 265542 -6106
rect 264986 -6662 265222 -6426
rect 265306 -6662 265542 -6426
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 289826 111218 290062 111454
rect 290146 111218 290382 111454
rect 289826 110898 290062 111134
rect 290146 110898 290382 111134
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 293546 150938 293782 151174
rect 293866 150938 294102 151174
rect 293546 150618 293782 150854
rect 293866 150618 294102 150854
rect 293546 114938 293782 115174
rect 293866 114938 294102 115174
rect 293546 114618 293782 114854
rect 293866 114618 294102 114854
rect 293546 78938 293782 79174
rect 293866 78938 294102 79174
rect 293546 78618 293782 78854
rect 293866 78618 294102 78854
rect 293546 42938 293782 43174
rect 293866 42938 294102 43174
rect 293546 42618 293782 42854
rect 293866 42618 294102 42854
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 293546 -2502 293782 -2266
rect 293866 -2502 294102 -2266
rect 293546 -2822 293782 -2586
rect 293866 -2822 294102 -2586
rect 297266 154658 297502 154894
rect 297586 154658 297822 154894
rect 297266 154338 297502 154574
rect 297586 154338 297822 154574
rect 297266 118658 297502 118894
rect 297586 118658 297822 118894
rect 297266 118338 297502 118574
rect 297586 118338 297822 118574
rect 297266 82658 297502 82894
rect 297586 82658 297822 82894
rect 297266 82338 297502 82574
rect 297586 82338 297822 82574
rect 297266 46658 297502 46894
rect 297586 46658 297822 46894
rect 297266 46338 297502 46574
rect 297586 46338 297822 46574
rect 297266 10658 297502 10894
rect 297586 10658 297822 10894
rect 297266 10338 297502 10574
rect 297586 10338 297822 10574
rect 297266 -4422 297502 -4186
rect 297586 -4422 297822 -4186
rect 297266 -4742 297502 -4506
rect 297586 -4742 297822 -4506
rect 300986 158378 301222 158614
rect 301306 158378 301542 158614
rect 300986 158058 301222 158294
rect 301306 158058 301542 158294
rect 300986 122378 301222 122614
rect 301306 122378 301542 122614
rect 300986 122058 301222 122294
rect 301306 122058 301542 122294
rect 300986 86378 301222 86614
rect 301306 86378 301542 86614
rect 300986 86058 301222 86294
rect 301306 86058 301542 86294
rect 300986 50378 301222 50614
rect 301306 50378 301542 50614
rect 300986 50058 301222 50294
rect 301306 50058 301542 50294
rect 300986 14378 301222 14614
rect 301306 14378 301542 14614
rect 300986 14058 301222 14294
rect 301306 14058 301542 14294
rect 282986 -7302 283222 -7066
rect 283306 -7302 283542 -7066
rect 282986 -7622 283222 -7386
rect 283306 -7622 283542 -7386
rect 307826 165218 308062 165454
rect 308146 165218 308382 165454
rect 307826 164898 308062 165134
rect 308146 164898 308382 165134
rect 307826 129218 308062 129454
rect 308146 129218 308382 129454
rect 307826 128898 308062 129134
rect 308146 128898 308382 129134
rect 307826 93218 308062 93454
rect 308146 93218 308382 93454
rect 307826 92898 308062 93134
rect 308146 92898 308382 93134
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -1542 308062 -1306
rect 308146 -1542 308382 -1306
rect 307826 -1862 308062 -1626
rect 308146 -1862 308382 -1626
rect 311546 168938 311782 169174
rect 311866 168938 312102 169174
rect 311546 168618 311782 168854
rect 311866 168618 312102 168854
rect 311546 132938 311782 133174
rect 311866 132938 312102 133174
rect 311546 132618 311782 132854
rect 311866 132618 312102 132854
rect 311546 96938 311782 97174
rect 311866 96938 312102 97174
rect 311546 96618 311782 96854
rect 311866 96618 312102 96854
rect 311546 60938 311782 61174
rect 311866 60938 312102 61174
rect 311546 60618 311782 60854
rect 311866 60618 312102 60854
rect 311546 24938 311782 25174
rect 311866 24938 312102 25174
rect 311546 24618 311782 24854
rect 311866 24618 312102 24854
rect 311546 -3462 311782 -3226
rect 311866 -3462 312102 -3226
rect 311546 -3782 311782 -3546
rect 311866 -3782 312102 -3546
rect 315266 172658 315502 172894
rect 315586 172658 315822 172894
rect 315266 172338 315502 172574
rect 315586 172338 315822 172574
rect 315266 136658 315502 136894
rect 315586 136658 315822 136894
rect 315266 136338 315502 136574
rect 315586 136338 315822 136574
rect 315266 100658 315502 100894
rect 315586 100658 315822 100894
rect 315266 100338 315502 100574
rect 315586 100338 315822 100574
rect 315266 64658 315502 64894
rect 315586 64658 315822 64894
rect 315266 64338 315502 64574
rect 315586 64338 315822 64574
rect 315266 28658 315502 28894
rect 315586 28658 315822 28894
rect 315266 28338 315502 28574
rect 315586 28338 315822 28574
rect 315266 -5382 315502 -5146
rect 315586 -5382 315822 -5146
rect 315266 -5702 315502 -5466
rect 315586 -5702 315822 -5466
rect 318986 176378 319222 176614
rect 319306 176378 319542 176614
rect 318986 176058 319222 176294
rect 319306 176058 319542 176294
rect 318986 140378 319222 140614
rect 319306 140378 319542 140614
rect 318986 140058 319222 140294
rect 319306 140058 319542 140294
rect 318986 104378 319222 104614
rect 319306 104378 319542 104614
rect 318986 104058 319222 104294
rect 319306 104058 319542 104294
rect 318986 68378 319222 68614
rect 319306 68378 319542 68614
rect 318986 68058 319222 68294
rect 319306 68058 319542 68294
rect 318986 32378 319222 32614
rect 319306 32378 319542 32614
rect 318986 32058 319222 32294
rect 319306 32058 319542 32294
rect 300986 -6342 301222 -6106
rect 301306 -6342 301542 -6106
rect 300986 -6662 301222 -6426
rect 301306 -6662 301542 -6426
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 325826 111218 326062 111454
rect 326146 111218 326382 111454
rect 325826 110898 326062 111134
rect 326146 110898 326382 111134
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 150938 329782 151174
rect 329866 150938 330102 151174
rect 329546 150618 329782 150854
rect 329866 150618 330102 150854
rect 329546 114938 329782 115174
rect 329866 114938 330102 115174
rect 329546 114618 329782 114854
rect 329866 114618 330102 114854
rect 329546 78938 329782 79174
rect 329866 78938 330102 79174
rect 329546 78618 329782 78854
rect 329866 78618 330102 78854
rect 329546 42938 329782 43174
rect 329866 42938 330102 43174
rect 329546 42618 329782 42854
rect 329866 42618 330102 42854
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 329546 -2502 329782 -2266
rect 329866 -2502 330102 -2266
rect 329546 -2822 329782 -2586
rect 329866 -2822 330102 -2586
rect 333266 154658 333502 154894
rect 333586 154658 333822 154894
rect 333266 154338 333502 154574
rect 333586 154338 333822 154574
rect 333266 118658 333502 118894
rect 333586 118658 333822 118894
rect 333266 118338 333502 118574
rect 333586 118338 333822 118574
rect 333266 82658 333502 82894
rect 333586 82658 333822 82894
rect 333266 82338 333502 82574
rect 333586 82338 333822 82574
rect 333266 46658 333502 46894
rect 333586 46658 333822 46894
rect 333266 46338 333502 46574
rect 333586 46338 333822 46574
rect 333266 10658 333502 10894
rect 333586 10658 333822 10894
rect 333266 10338 333502 10574
rect 333586 10338 333822 10574
rect 333266 -4422 333502 -4186
rect 333586 -4422 333822 -4186
rect 333266 -4742 333502 -4506
rect 333586 -4742 333822 -4506
rect 336986 158378 337222 158614
rect 337306 158378 337542 158614
rect 336986 158058 337222 158294
rect 337306 158058 337542 158294
rect 336986 122378 337222 122614
rect 337306 122378 337542 122614
rect 336986 122058 337222 122294
rect 337306 122058 337542 122294
rect 336986 86378 337222 86614
rect 337306 86378 337542 86614
rect 336986 86058 337222 86294
rect 337306 86058 337542 86294
rect 336986 50378 337222 50614
rect 337306 50378 337542 50614
rect 336986 50058 337222 50294
rect 337306 50058 337542 50294
rect 336986 14378 337222 14614
rect 337306 14378 337542 14614
rect 336986 14058 337222 14294
rect 337306 14058 337542 14294
rect 318986 -7302 319222 -7066
rect 319306 -7302 319542 -7066
rect 318986 -7622 319222 -7386
rect 319306 -7622 319542 -7386
rect 343826 165218 344062 165454
rect 344146 165218 344382 165454
rect 343826 164898 344062 165134
rect 344146 164898 344382 165134
rect 343826 129218 344062 129454
rect 344146 129218 344382 129454
rect 343826 128898 344062 129134
rect 344146 128898 344382 129134
rect 343826 93218 344062 93454
rect 344146 93218 344382 93454
rect 343826 92898 344062 93134
rect 344146 92898 344382 93134
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -1542 344062 -1306
rect 344146 -1542 344382 -1306
rect 343826 -1862 344062 -1626
rect 344146 -1862 344382 -1626
rect 347546 168938 347782 169174
rect 347866 168938 348102 169174
rect 347546 168618 347782 168854
rect 347866 168618 348102 168854
rect 347546 132938 347782 133174
rect 347866 132938 348102 133174
rect 347546 132618 347782 132854
rect 347866 132618 348102 132854
rect 347546 96938 347782 97174
rect 347866 96938 348102 97174
rect 347546 96618 347782 96854
rect 347866 96618 348102 96854
rect 347546 60938 347782 61174
rect 347866 60938 348102 61174
rect 347546 60618 347782 60854
rect 347866 60618 348102 60854
rect 347546 24938 347782 25174
rect 347866 24938 348102 25174
rect 347546 24618 347782 24854
rect 347866 24618 348102 24854
rect 347546 -3462 347782 -3226
rect 347866 -3462 348102 -3226
rect 347546 -3782 347782 -3546
rect 347866 -3782 348102 -3546
rect 351266 172658 351502 172894
rect 351586 172658 351822 172894
rect 351266 172338 351502 172574
rect 351586 172338 351822 172574
rect 351266 136658 351502 136894
rect 351586 136658 351822 136894
rect 351266 136338 351502 136574
rect 351586 136338 351822 136574
rect 351266 100658 351502 100894
rect 351586 100658 351822 100894
rect 351266 100338 351502 100574
rect 351586 100338 351822 100574
rect 351266 64658 351502 64894
rect 351586 64658 351822 64894
rect 351266 64338 351502 64574
rect 351586 64338 351822 64574
rect 351266 28658 351502 28894
rect 351586 28658 351822 28894
rect 351266 28338 351502 28574
rect 351586 28338 351822 28574
rect 351266 -5382 351502 -5146
rect 351586 -5382 351822 -5146
rect 351266 -5702 351502 -5466
rect 351586 -5702 351822 -5466
rect 354986 176378 355222 176614
rect 355306 176378 355542 176614
rect 354986 176058 355222 176294
rect 355306 176058 355542 176294
rect 354986 140378 355222 140614
rect 355306 140378 355542 140614
rect 354986 140058 355222 140294
rect 355306 140058 355542 140294
rect 354986 104378 355222 104614
rect 355306 104378 355542 104614
rect 354986 104058 355222 104294
rect 355306 104058 355542 104294
rect 354986 68378 355222 68614
rect 355306 68378 355542 68614
rect 354986 68058 355222 68294
rect 355306 68058 355542 68294
rect 354986 32378 355222 32614
rect 355306 32378 355542 32614
rect 354986 32058 355222 32294
rect 355306 32058 355542 32294
rect 336986 -6342 337222 -6106
rect 337306 -6342 337542 -6106
rect 336986 -6662 337222 -6426
rect 337306 -6662 337542 -6426
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 365546 150938 365782 151174
rect 365866 150938 366102 151174
rect 365546 150618 365782 150854
rect 365866 150618 366102 150854
rect 365546 114938 365782 115174
rect 365866 114938 366102 115174
rect 365546 114618 365782 114854
rect 365866 114618 366102 114854
rect 365546 78938 365782 79174
rect 365866 78938 366102 79174
rect 365546 78618 365782 78854
rect 365866 78618 366102 78854
rect 365546 42938 365782 43174
rect 365866 42938 366102 43174
rect 365546 42618 365782 42854
rect 365866 42618 366102 42854
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 365546 -2502 365782 -2266
rect 365866 -2502 366102 -2266
rect 365546 -2822 365782 -2586
rect 365866 -2822 366102 -2586
rect 369266 154658 369502 154894
rect 369586 154658 369822 154894
rect 369266 154338 369502 154574
rect 369586 154338 369822 154574
rect 369266 118658 369502 118894
rect 369586 118658 369822 118894
rect 369266 118338 369502 118574
rect 369586 118338 369822 118574
rect 369266 82658 369502 82894
rect 369586 82658 369822 82894
rect 369266 82338 369502 82574
rect 369586 82338 369822 82574
rect 369266 46658 369502 46894
rect 369586 46658 369822 46894
rect 369266 46338 369502 46574
rect 369586 46338 369822 46574
rect 369266 10658 369502 10894
rect 369586 10658 369822 10894
rect 369266 10338 369502 10574
rect 369586 10338 369822 10574
rect 369266 -4422 369502 -4186
rect 369586 -4422 369822 -4186
rect 369266 -4742 369502 -4506
rect 369586 -4742 369822 -4506
rect 372986 158378 373222 158614
rect 373306 158378 373542 158614
rect 372986 158058 373222 158294
rect 373306 158058 373542 158294
rect 372986 122378 373222 122614
rect 373306 122378 373542 122614
rect 372986 122058 373222 122294
rect 373306 122058 373542 122294
rect 372986 86378 373222 86614
rect 373306 86378 373542 86614
rect 372986 86058 373222 86294
rect 373306 86058 373542 86294
rect 372986 50378 373222 50614
rect 373306 50378 373542 50614
rect 372986 50058 373222 50294
rect 373306 50058 373542 50294
rect 372986 14378 373222 14614
rect 373306 14378 373542 14614
rect 372986 14058 373222 14294
rect 373306 14058 373542 14294
rect 354986 -7302 355222 -7066
rect 355306 -7302 355542 -7066
rect 354986 -7622 355222 -7386
rect 355306 -7622 355542 -7386
rect 379826 165218 380062 165454
rect 380146 165218 380382 165454
rect 379826 164898 380062 165134
rect 380146 164898 380382 165134
rect 379826 129218 380062 129454
rect 380146 129218 380382 129454
rect 379826 128898 380062 129134
rect 380146 128898 380382 129134
rect 379826 93218 380062 93454
rect 380146 93218 380382 93454
rect 379826 92898 380062 93134
rect 380146 92898 380382 93134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -1542 380062 -1306
rect 380146 -1542 380382 -1306
rect 379826 -1862 380062 -1626
rect 380146 -1862 380382 -1626
rect 383546 168938 383782 169174
rect 383866 168938 384102 169174
rect 383546 168618 383782 168854
rect 383866 168618 384102 168854
rect 383546 132938 383782 133174
rect 383866 132938 384102 133174
rect 383546 132618 383782 132854
rect 383866 132618 384102 132854
rect 383546 96938 383782 97174
rect 383866 96938 384102 97174
rect 383546 96618 383782 96854
rect 383866 96618 384102 96854
rect 383546 60938 383782 61174
rect 383866 60938 384102 61174
rect 383546 60618 383782 60854
rect 383866 60618 384102 60854
rect 383546 24938 383782 25174
rect 383866 24938 384102 25174
rect 383546 24618 383782 24854
rect 383866 24618 384102 24854
rect 383546 -3462 383782 -3226
rect 383866 -3462 384102 -3226
rect 383546 -3782 383782 -3546
rect 383866 -3782 384102 -3546
rect 387266 172658 387502 172894
rect 387586 172658 387822 172894
rect 387266 172338 387502 172574
rect 387586 172338 387822 172574
rect 387266 136658 387502 136894
rect 387586 136658 387822 136894
rect 387266 136338 387502 136574
rect 387586 136338 387822 136574
rect 387266 100658 387502 100894
rect 387586 100658 387822 100894
rect 387266 100338 387502 100574
rect 387586 100338 387822 100574
rect 387266 64658 387502 64894
rect 387586 64658 387822 64894
rect 387266 64338 387502 64574
rect 387586 64338 387822 64574
rect 387266 28658 387502 28894
rect 387586 28658 387822 28894
rect 387266 28338 387502 28574
rect 387586 28338 387822 28574
rect 387266 -5382 387502 -5146
rect 387586 -5382 387822 -5146
rect 387266 -5702 387502 -5466
rect 387586 -5702 387822 -5466
rect 390986 176378 391222 176614
rect 391306 176378 391542 176614
rect 390986 176058 391222 176294
rect 391306 176058 391542 176294
rect 390986 140378 391222 140614
rect 391306 140378 391542 140614
rect 390986 140058 391222 140294
rect 391306 140058 391542 140294
rect 390986 104378 391222 104614
rect 391306 104378 391542 104614
rect 390986 104058 391222 104294
rect 391306 104058 391542 104294
rect 390986 68378 391222 68614
rect 391306 68378 391542 68614
rect 390986 68058 391222 68294
rect 391306 68058 391542 68294
rect 390986 32378 391222 32614
rect 391306 32378 391542 32614
rect 390986 32058 391222 32294
rect 391306 32058 391542 32294
rect 372986 -6342 373222 -6106
rect 373306 -6342 373542 -6106
rect 372986 -6662 373222 -6426
rect 373306 -6662 373542 -6426
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 150938 401782 151174
rect 401866 150938 402102 151174
rect 401546 150618 401782 150854
rect 401866 150618 402102 150854
rect 401546 114938 401782 115174
rect 401866 114938 402102 115174
rect 401546 114618 401782 114854
rect 401866 114618 402102 114854
rect 401546 78938 401782 79174
rect 401866 78938 402102 79174
rect 401546 78618 401782 78854
rect 401866 78618 402102 78854
rect 401546 42938 401782 43174
rect 401866 42938 402102 43174
rect 401546 42618 401782 42854
rect 401866 42618 402102 42854
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -2502 401782 -2266
rect 401866 -2502 402102 -2266
rect 401546 -2822 401782 -2586
rect 401866 -2822 402102 -2586
rect 405266 154658 405502 154894
rect 405586 154658 405822 154894
rect 405266 154338 405502 154574
rect 405586 154338 405822 154574
rect 405266 118658 405502 118894
rect 405586 118658 405822 118894
rect 405266 118338 405502 118574
rect 405586 118338 405822 118574
rect 405266 82658 405502 82894
rect 405586 82658 405822 82894
rect 405266 82338 405502 82574
rect 405586 82338 405822 82574
rect 405266 46658 405502 46894
rect 405586 46658 405822 46894
rect 405266 46338 405502 46574
rect 405586 46338 405822 46574
rect 405266 10658 405502 10894
rect 405586 10658 405822 10894
rect 405266 10338 405502 10574
rect 405586 10338 405822 10574
rect 405266 -4422 405502 -4186
rect 405586 -4422 405822 -4186
rect 405266 -4742 405502 -4506
rect 405586 -4742 405822 -4506
rect 408986 158378 409222 158614
rect 409306 158378 409542 158614
rect 408986 158058 409222 158294
rect 409306 158058 409542 158294
rect 408986 122378 409222 122614
rect 409306 122378 409542 122614
rect 408986 122058 409222 122294
rect 409306 122058 409542 122294
rect 408986 86378 409222 86614
rect 409306 86378 409542 86614
rect 408986 86058 409222 86294
rect 409306 86058 409542 86294
rect 408986 50378 409222 50614
rect 409306 50378 409542 50614
rect 408986 50058 409222 50294
rect 409306 50058 409542 50294
rect 408986 14378 409222 14614
rect 409306 14378 409542 14614
rect 408986 14058 409222 14294
rect 409306 14058 409542 14294
rect 390986 -7302 391222 -7066
rect 391306 -7302 391542 -7066
rect 390986 -7622 391222 -7386
rect 391306 -7622 391542 -7386
rect 415826 165218 416062 165454
rect 416146 165218 416382 165454
rect 415826 164898 416062 165134
rect 416146 164898 416382 165134
rect 415826 129218 416062 129454
rect 416146 129218 416382 129454
rect 415826 128898 416062 129134
rect 416146 128898 416382 129134
rect 415826 93218 416062 93454
rect 416146 93218 416382 93454
rect 415826 92898 416062 93134
rect 416146 92898 416382 93134
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -1542 416062 -1306
rect 416146 -1542 416382 -1306
rect 415826 -1862 416062 -1626
rect 416146 -1862 416382 -1626
rect 419546 168938 419782 169174
rect 419866 168938 420102 169174
rect 419546 168618 419782 168854
rect 419866 168618 420102 168854
rect 419546 132938 419782 133174
rect 419866 132938 420102 133174
rect 419546 132618 419782 132854
rect 419866 132618 420102 132854
rect 419546 96938 419782 97174
rect 419866 96938 420102 97174
rect 419546 96618 419782 96854
rect 419866 96618 420102 96854
rect 419546 60938 419782 61174
rect 419866 60938 420102 61174
rect 419546 60618 419782 60854
rect 419866 60618 420102 60854
rect 419546 24938 419782 25174
rect 419866 24938 420102 25174
rect 419546 24618 419782 24854
rect 419866 24618 420102 24854
rect 419546 -3462 419782 -3226
rect 419866 -3462 420102 -3226
rect 419546 -3782 419782 -3546
rect 419866 -3782 420102 -3546
rect 423266 172658 423502 172894
rect 423586 172658 423822 172894
rect 423266 172338 423502 172574
rect 423586 172338 423822 172574
rect 423266 136658 423502 136894
rect 423586 136658 423822 136894
rect 423266 136338 423502 136574
rect 423586 136338 423822 136574
rect 423266 100658 423502 100894
rect 423586 100658 423822 100894
rect 423266 100338 423502 100574
rect 423586 100338 423822 100574
rect 423266 64658 423502 64894
rect 423586 64658 423822 64894
rect 423266 64338 423502 64574
rect 423586 64338 423822 64574
rect 423266 28658 423502 28894
rect 423586 28658 423822 28894
rect 423266 28338 423502 28574
rect 423586 28338 423822 28574
rect 423266 -5382 423502 -5146
rect 423586 -5382 423822 -5146
rect 423266 -5702 423502 -5466
rect 423586 -5702 423822 -5466
rect 426986 176378 427222 176614
rect 427306 176378 427542 176614
rect 426986 176058 427222 176294
rect 427306 176058 427542 176294
rect 426986 140378 427222 140614
rect 427306 140378 427542 140614
rect 426986 140058 427222 140294
rect 427306 140058 427542 140294
rect 426986 104378 427222 104614
rect 427306 104378 427542 104614
rect 426986 104058 427222 104294
rect 427306 104058 427542 104294
rect 426986 68378 427222 68614
rect 427306 68378 427542 68614
rect 426986 68058 427222 68294
rect 427306 68058 427542 68294
rect 426986 32378 427222 32614
rect 427306 32378 427542 32614
rect 426986 32058 427222 32294
rect 427306 32058 427542 32294
rect 408986 -6342 409222 -6106
rect 409306 -6342 409542 -6106
rect 408986 -6662 409222 -6426
rect 409306 -6662 409542 -6426
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 150938 437782 151174
rect 437866 150938 438102 151174
rect 437546 150618 437782 150854
rect 437866 150618 438102 150854
rect 437546 114938 437782 115174
rect 437866 114938 438102 115174
rect 437546 114618 437782 114854
rect 437866 114618 438102 114854
rect 437546 78938 437782 79174
rect 437866 78938 438102 79174
rect 437546 78618 437782 78854
rect 437866 78618 438102 78854
rect 437546 42938 437782 43174
rect 437866 42938 438102 43174
rect 437546 42618 437782 42854
rect 437866 42618 438102 42854
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 437546 -2502 437782 -2266
rect 437866 -2502 438102 -2266
rect 437546 -2822 437782 -2586
rect 437866 -2822 438102 -2586
rect 441266 154658 441502 154894
rect 441586 154658 441822 154894
rect 441266 154338 441502 154574
rect 441586 154338 441822 154574
rect 441266 118658 441502 118894
rect 441586 118658 441822 118894
rect 441266 118338 441502 118574
rect 441586 118338 441822 118574
rect 441266 82658 441502 82894
rect 441586 82658 441822 82894
rect 441266 82338 441502 82574
rect 441586 82338 441822 82574
rect 441266 46658 441502 46894
rect 441586 46658 441822 46894
rect 441266 46338 441502 46574
rect 441586 46338 441822 46574
rect 441266 10658 441502 10894
rect 441586 10658 441822 10894
rect 441266 10338 441502 10574
rect 441586 10338 441822 10574
rect 441266 -4422 441502 -4186
rect 441586 -4422 441822 -4186
rect 441266 -4742 441502 -4506
rect 441586 -4742 441822 -4506
rect 444986 158378 445222 158614
rect 445306 158378 445542 158614
rect 444986 158058 445222 158294
rect 445306 158058 445542 158294
rect 444986 122378 445222 122614
rect 445306 122378 445542 122614
rect 444986 122058 445222 122294
rect 445306 122058 445542 122294
rect 444986 86378 445222 86614
rect 445306 86378 445542 86614
rect 444986 86058 445222 86294
rect 445306 86058 445542 86294
rect 444986 50378 445222 50614
rect 445306 50378 445542 50614
rect 444986 50058 445222 50294
rect 445306 50058 445542 50294
rect 444986 14378 445222 14614
rect 445306 14378 445542 14614
rect 444986 14058 445222 14294
rect 445306 14058 445542 14294
rect 426986 -7302 427222 -7066
rect 427306 -7302 427542 -7066
rect 426986 -7622 427222 -7386
rect 427306 -7622 427542 -7386
rect 451826 165218 452062 165454
rect 452146 165218 452382 165454
rect 451826 164898 452062 165134
rect 452146 164898 452382 165134
rect 451826 129218 452062 129454
rect 452146 129218 452382 129454
rect 451826 128898 452062 129134
rect 452146 128898 452382 129134
rect 451826 93218 452062 93454
rect 452146 93218 452382 93454
rect 451826 92898 452062 93134
rect 452146 92898 452382 93134
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -1542 452062 -1306
rect 452146 -1542 452382 -1306
rect 451826 -1862 452062 -1626
rect 452146 -1862 452382 -1626
rect 455546 168938 455782 169174
rect 455866 168938 456102 169174
rect 455546 168618 455782 168854
rect 455866 168618 456102 168854
rect 455546 132938 455782 133174
rect 455866 132938 456102 133174
rect 455546 132618 455782 132854
rect 455866 132618 456102 132854
rect 455546 96938 455782 97174
rect 455866 96938 456102 97174
rect 455546 96618 455782 96854
rect 455866 96618 456102 96854
rect 455546 60938 455782 61174
rect 455866 60938 456102 61174
rect 455546 60618 455782 60854
rect 455866 60618 456102 60854
rect 455546 24938 455782 25174
rect 455866 24938 456102 25174
rect 455546 24618 455782 24854
rect 455866 24618 456102 24854
rect 455546 -3462 455782 -3226
rect 455866 -3462 456102 -3226
rect 455546 -3782 455782 -3546
rect 455866 -3782 456102 -3546
rect 459266 172658 459502 172894
rect 459586 172658 459822 172894
rect 459266 172338 459502 172574
rect 459586 172338 459822 172574
rect 459266 136658 459502 136894
rect 459586 136658 459822 136894
rect 459266 136338 459502 136574
rect 459586 136338 459822 136574
rect 459266 100658 459502 100894
rect 459586 100658 459822 100894
rect 459266 100338 459502 100574
rect 459586 100338 459822 100574
rect 459266 64658 459502 64894
rect 459586 64658 459822 64894
rect 459266 64338 459502 64574
rect 459586 64338 459822 64574
rect 459266 28658 459502 28894
rect 459586 28658 459822 28894
rect 459266 28338 459502 28574
rect 459586 28338 459822 28574
rect 459266 -5382 459502 -5146
rect 459586 -5382 459822 -5146
rect 459266 -5702 459502 -5466
rect 459586 -5702 459822 -5466
rect 462986 176378 463222 176614
rect 463306 176378 463542 176614
rect 462986 176058 463222 176294
rect 463306 176058 463542 176294
rect 462986 140378 463222 140614
rect 463306 140378 463542 140614
rect 462986 140058 463222 140294
rect 463306 140058 463542 140294
rect 462986 104378 463222 104614
rect 463306 104378 463542 104614
rect 462986 104058 463222 104294
rect 463306 104058 463542 104294
rect 462986 68378 463222 68614
rect 463306 68378 463542 68614
rect 462986 68058 463222 68294
rect 463306 68058 463542 68294
rect 462986 32378 463222 32614
rect 463306 32378 463542 32614
rect 462986 32058 463222 32294
rect 463306 32058 463542 32294
rect 444986 -6342 445222 -6106
rect 445306 -6342 445542 -6106
rect 444986 -6662 445222 -6426
rect 445306 -6662 445542 -6426
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 150938 473782 151174
rect 473866 150938 474102 151174
rect 473546 150618 473782 150854
rect 473866 150618 474102 150854
rect 473546 114938 473782 115174
rect 473866 114938 474102 115174
rect 473546 114618 473782 114854
rect 473866 114618 474102 114854
rect 473546 78938 473782 79174
rect 473866 78938 474102 79174
rect 473546 78618 473782 78854
rect 473866 78618 474102 78854
rect 473546 42938 473782 43174
rect 473866 42938 474102 43174
rect 473546 42618 473782 42854
rect 473866 42618 474102 42854
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -2502 473782 -2266
rect 473866 -2502 474102 -2266
rect 473546 -2822 473782 -2586
rect 473866 -2822 474102 -2586
rect 477266 154658 477502 154894
rect 477586 154658 477822 154894
rect 477266 154338 477502 154574
rect 477586 154338 477822 154574
rect 477266 118658 477502 118894
rect 477586 118658 477822 118894
rect 477266 118338 477502 118574
rect 477586 118338 477822 118574
rect 477266 82658 477502 82894
rect 477586 82658 477822 82894
rect 477266 82338 477502 82574
rect 477586 82338 477822 82574
rect 477266 46658 477502 46894
rect 477586 46658 477822 46894
rect 477266 46338 477502 46574
rect 477586 46338 477822 46574
rect 477266 10658 477502 10894
rect 477586 10658 477822 10894
rect 477266 10338 477502 10574
rect 477586 10338 477822 10574
rect 477266 -4422 477502 -4186
rect 477586 -4422 477822 -4186
rect 477266 -4742 477502 -4506
rect 477586 -4742 477822 -4506
rect 480986 158378 481222 158614
rect 481306 158378 481542 158614
rect 480986 158058 481222 158294
rect 481306 158058 481542 158294
rect 480986 122378 481222 122614
rect 481306 122378 481542 122614
rect 480986 122058 481222 122294
rect 481306 122058 481542 122294
rect 480986 86378 481222 86614
rect 481306 86378 481542 86614
rect 480986 86058 481222 86294
rect 481306 86058 481542 86294
rect 480986 50378 481222 50614
rect 481306 50378 481542 50614
rect 480986 50058 481222 50294
rect 481306 50058 481542 50294
rect 480986 14378 481222 14614
rect 481306 14378 481542 14614
rect 480986 14058 481222 14294
rect 481306 14058 481542 14294
rect 462986 -7302 463222 -7066
rect 463306 -7302 463542 -7066
rect 462986 -7622 463222 -7386
rect 463306 -7622 463542 -7386
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 487826 129218 488062 129454
rect 488146 129218 488382 129454
rect 487826 128898 488062 129134
rect 488146 128898 488382 129134
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -1542 488062 -1306
rect 488146 -1542 488382 -1306
rect 487826 -1862 488062 -1626
rect 488146 -1862 488382 -1626
rect 491546 168938 491782 169174
rect 491866 168938 492102 169174
rect 491546 168618 491782 168854
rect 491866 168618 492102 168854
rect 491546 132938 491782 133174
rect 491866 132938 492102 133174
rect 491546 132618 491782 132854
rect 491866 132618 492102 132854
rect 491546 96938 491782 97174
rect 491866 96938 492102 97174
rect 491546 96618 491782 96854
rect 491866 96618 492102 96854
rect 491546 60938 491782 61174
rect 491866 60938 492102 61174
rect 491546 60618 491782 60854
rect 491866 60618 492102 60854
rect 491546 24938 491782 25174
rect 491866 24938 492102 25174
rect 491546 24618 491782 24854
rect 491866 24618 492102 24854
rect 491546 -3462 491782 -3226
rect 491866 -3462 492102 -3226
rect 491546 -3782 491782 -3546
rect 491866 -3782 492102 -3546
rect 495266 172658 495502 172894
rect 495586 172658 495822 172894
rect 495266 172338 495502 172574
rect 495586 172338 495822 172574
rect 495266 136658 495502 136894
rect 495586 136658 495822 136894
rect 495266 136338 495502 136574
rect 495586 136338 495822 136574
rect 495266 100658 495502 100894
rect 495586 100658 495822 100894
rect 495266 100338 495502 100574
rect 495586 100338 495822 100574
rect 495266 64658 495502 64894
rect 495586 64658 495822 64894
rect 495266 64338 495502 64574
rect 495586 64338 495822 64574
rect 495266 28658 495502 28894
rect 495586 28658 495822 28894
rect 495266 28338 495502 28574
rect 495586 28338 495822 28574
rect 495266 -5382 495502 -5146
rect 495586 -5382 495822 -5146
rect 495266 -5702 495502 -5466
rect 495586 -5702 495822 -5466
rect 498986 176378 499222 176614
rect 499306 176378 499542 176614
rect 498986 176058 499222 176294
rect 499306 176058 499542 176294
rect 498986 140378 499222 140614
rect 499306 140378 499542 140614
rect 498986 140058 499222 140294
rect 499306 140058 499542 140294
rect 498986 104378 499222 104614
rect 499306 104378 499542 104614
rect 498986 104058 499222 104294
rect 499306 104058 499542 104294
rect 498986 68378 499222 68614
rect 499306 68378 499542 68614
rect 498986 68058 499222 68294
rect 499306 68058 499542 68294
rect 498986 32378 499222 32614
rect 499306 32378 499542 32614
rect 498986 32058 499222 32294
rect 499306 32058 499542 32294
rect 480986 -6342 481222 -6106
rect 481306 -6342 481542 -6106
rect 480986 -6662 481222 -6426
rect 481306 -6662 481542 -6426
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 690938 509782 691174
rect 509866 690938 510102 691174
rect 509546 690618 509782 690854
rect 509866 690618 510102 690854
rect 509546 654938 509782 655174
rect 509866 654938 510102 655174
rect 509546 654618 509782 654854
rect 509866 654618 510102 654854
rect 509546 618938 509782 619174
rect 509866 618938 510102 619174
rect 509546 618618 509782 618854
rect 509866 618618 510102 618854
rect 509546 582938 509782 583174
rect 509866 582938 510102 583174
rect 509546 582618 509782 582854
rect 509866 582618 510102 582854
rect 509546 546938 509782 547174
rect 509866 546938 510102 547174
rect 509546 546618 509782 546854
rect 509866 546618 510102 546854
rect 509546 510938 509782 511174
rect 509866 510938 510102 511174
rect 509546 510618 509782 510854
rect 509866 510618 510102 510854
rect 509546 474938 509782 475174
rect 509866 474938 510102 475174
rect 509546 474618 509782 474854
rect 509866 474618 510102 474854
rect 509546 438938 509782 439174
rect 509866 438938 510102 439174
rect 509546 438618 509782 438854
rect 509866 438618 510102 438854
rect 509546 402938 509782 403174
rect 509866 402938 510102 403174
rect 509546 402618 509782 402854
rect 509866 402618 510102 402854
rect 509546 366938 509782 367174
rect 509866 366938 510102 367174
rect 509546 366618 509782 366854
rect 509866 366618 510102 366854
rect 509546 330938 509782 331174
rect 509866 330938 510102 331174
rect 509546 330618 509782 330854
rect 509866 330618 510102 330854
rect 509546 294938 509782 295174
rect 509866 294938 510102 295174
rect 509546 294618 509782 294854
rect 509866 294618 510102 294854
rect 509546 258938 509782 259174
rect 509866 258938 510102 259174
rect 509546 258618 509782 258854
rect 509866 258618 510102 258854
rect 509546 222938 509782 223174
rect 509866 222938 510102 223174
rect 509546 222618 509782 222854
rect 509866 222618 510102 222854
rect 509546 186938 509782 187174
rect 509866 186938 510102 187174
rect 509546 186618 509782 186854
rect 509866 186618 510102 186854
rect 509546 150938 509782 151174
rect 509866 150938 510102 151174
rect 509546 150618 509782 150854
rect 509866 150618 510102 150854
rect 509546 114938 509782 115174
rect 509866 114938 510102 115174
rect 509546 114618 509782 114854
rect 509866 114618 510102 114854
rect 509546 78938 509782 79174
rect 509866 78938 510102 79174
rect 509546 78618 509782 78854
rect 509866 78618 510102 78854
rect 509546 42938 509782 43174
rect 509866 42938 510102 43174
rect 509546 42618 509782 42854
rect 509866 42618 510102 42854
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -2502 509782 -2266
rect 509866 -2502 510102 -2266
rect 509546 -2822 509782 -2586
rect 509866 -2822 510102 -2586
rect 513266 694658 513502 694894
rect 513586 694658 513822 694894
rect 513266 694338 513502 694574
rect 513586 694338 513822 694574
rect 513266 658658 513502 658894
rect 513586 658658 513822 658894
rect 513266 658338 513502 658574
rect 513586 658338 513822 658574
rect 513266 622658 513502 622894
rect 513586 622658 513822 622894
rect 513266 622338 513502 622574
rect 513586 622338 513822 622574
rect 513266 586658 513502 586894
rect 513586 586658 513822 586894
rect 513266 586338 513502 586574
rect 513586 586338 513822 586574
rect 513266 550658 513502 550894
rect 513586 550658 513822 550894
rect 513266 550338 513502 550574
rect 513586 550338 513822 550574
rect 513266 514658 513502 514894
rect 513586 514658 513822 514894
rect 513266 514338 513502 514574
rect 513586 514338 513822 514574
rect 513266 478658 513502 478894
rect 513586 478658 513822 478894
rect 513266 478338 513502 478574
rect 513586 478338 513822 478574
rect 513266 442658 513502 442894
rect 513586 442658 513822 442894
rect 513266 442338 513502 442574
rect 513586 442338 513822 442574
rect 513266 406658 513502 406894
rect 513586 406658 513822 406894
rect 513266 406338 513502 406574
rect 513586 406338 513822 406574
rect 513266 370658 513502 370894
rect 513586 370658 513822 370894
rect 513266 370338 513502 370574
rect 513586 370338 513822 370574
rect 513266 334658 513502 334894
rect 513586 334658 513822 334894
rect 513266 334338 513502 334574
rect 513586 334338 513822 334574
rect 513266 298658 513502 298894
rect 513586 298658 513822 298894
rect 513266 298338 513502 298574
rect 513586 298338 513822 298574
rect 513266 262658 513502 262894
rect 513586 262658 513822 262894
rect 513266 262338 513502 262574
rect 513586 262338 513822 262574
rect 513266 226658 513502 226894
rect 513586 226658 513822 226894
rect 513266 226338 513502 226574
rect 513586 226338 513822 226574
rect 513266 190658 513502 190894
rect 513586 190658 513822 190894
rect 513266 190338 513502 190574
rect 513586 190338 513822 190574
rect 513266 154658 513502 154894
rect 513586 154658 513822 154894
rect 513266 154338 513502 154574
rect 513586 154338 513822 154574
rect 513266 118658 513502 118894
rect 513586 118658 513822 118894
rect 513266 118338 513502 118574
rect 513586 118338 513822 118574
rect 513266 82658 513502 82894
rect 513586 82658 513822 82894
rect 513266 82338 513502 82574
rect 513586 82338 513822 82574
rect 513266 46658 513502 46894
rect 513586 46658 513822 46894
rect 513266 46338 513502 46574
rect 513586 46338 513822 46574
rect 513266 10658 513502 10894
rect 513586 10658 513822 10894
rect 513266 10338 513502 10574
rect 513586 10338 513822 10574
rect 513266 -4422 513502 -4186
rect 513586 -4422 513822 -4186
rect 513266 -4742 513502 -4506
rect 513586 -4742 513822 -4506
rect 534986 711322 535222 711558
rect 535306 711322 535542 711558
rect 534986 711002 535222 711238
rect 535306 711002 535542 711238
rect 531266 709402 531502 709638
rect 531586 709402 531822 709638
rect 531266 709082 531502 709318
rect 531586 709082 531822 709318
rect 527546 707482 527782 707718
rect 527866 707482 528102 707718
rect 527546 707162 527782 707398
rect 527866 707162 528102 707398
rect 516986 698378 517222 698614
rect 517306 698378 517542 698614
rect 516986 698058 517222 698294
rect 517306 698058 517542 698294
rect 516986 662378 517222 662614
rect 517306 662378 517542 662614
rect 516986 662058 517222 662294
rect 517306 662058 517542 662294
rect 516986 626378 517222 626614
rect 517306 626378 517542 626614
rect 516986 626058 517222 626294
rect 517306 626058 517542 626294
rect 516986 590378 517222 590614
rect 517306 590378 517542 590614
rect 516986 590058 517222 590294
rect 517306 590058 517542 590294
rect 516986 554378 517222 554614
rect 517306 554378 517542 554614
rect 516986 554058 517222 554294
rect 517306 554058 517542 554294
rect 516986 518378 517222 518614
rect 517306 518378 517542 518614
rect 516986 518058 517222 518294
rect 517306 518058 517542 518294
rect 516986 482378 517222 482614
rect 517306 482378 517542 482614
rect 516986 482058 517222 482294
rect 517306 482058 517542 482294
rect 516986 446378 517222 446614
rect 517306 446378 517542 446614
rect 516986 446058 517222 446294
rect 517306 446058 517542 446294
rect 516986 410378 517222 410614
rect 517306 410378 517542 410614
rect 516986 410058 517222 410294
rect 517306 410058 517542 410294
rect 516986 374378 517222 374614
rect 517306 374378 517542 374614
rect 516986 374058 517222 374294
rect 517306 374058 517542 374294
rect 516986 338378 517222 338614
rect 517306 338378 517542 338614
rect 516986 338058 517222 338294
rect 517306 338058 517542 338294
rect 516986 302378 517222 302614
rect 517306 302378 517542 302614
rect 516986 302058 517222 302294
rect 517306 302058 517542 302294
rect 516986 266378 517222 266614
rect 517306 266378 517542 266614
rect 516986 266058 517222 266294
rect 517306 266058 517542 266294
rect 516986 230378 517222 230614
rect 517306 230378 517542 230614
rect 516986 230058 517222 230294
rect 517306 230058 517542 230294
rect 516986 194378 517222 194614
rect 517306 194378 517542 194614
rect 516986 194058 517222 194294
rect 517306 194058 517542 194294
rect 516986 158378 517222 158614
rect 517306 158378 517542 158614
rect 516986 158058 517222 158294
rect 517306 158058 517542 158294
rect 516986 122378 517222 122614
rect 517306 122378 517542 122614
rect 516986 122058 517222 122294
rect 517306 122058 517542 122294
rect 516986 86378 517222 86614
rect 517306 86378 517542 86614
rect 516986 86058 517222 86294
rect 517306 86058 517542 86294
rect 516986 50378 517222 50614
rect 517306 50378 517542 50614
rect 516986 50058 517222 50294
rect 517306 50058 517542 50294
rect 516986 14378 517222 14614
rect 517306 14378 517542 14614
rect 516986 14058 517222 14294
rect 517306 14058 517542 14294
rect 498986 -7302 499222 -7066
rect 499306 -7302 499542 -7066
rect 498986 -7622 499222 -7386
rect 499306 -7622 499542 -7386
rect 523826 705562 524062 705798
rect 524146 705562 524382 705798
rect 523826 705242 524062 705478
rect 524146 705242 524382 705478
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -1542 524062 -1306
rect 524146 -1542 524382 -1306
rect 523826 -1862 524062 -1626
rect 524146 -1862 524382 -1626
rect 527546 672938 527782 673174
rect 527866 672938 528102 673174
rect 527546 672618 527782 672854
rect 527866 672618 528102 672854
rect 527546 636938 527782 637174
rect 527866 636938 528102 637174
rect 527546 636618 527782 636854
rect 527866 636618 528102 636854
rect 527546 600938 527782 601174
rect 527866 600938 528102 601174
rect 527546 600618 527782 600854
rect 527866 600618 528102 600854
rect 527546 564938 527782 565174
rect 527866 564938 528102 565174
rect 527546 564618 527782 564854
rect 527866 564618 528102 564854
rect 527546 528938 527782 529174
rect 527866 528938 528102 529174
rect 527546 528618 527782 528854
rect 527866 528618 528102 528854
rect 527546 492938 527782 493174
rect 527866 492938 528102 493174
rect 527546 492618 527782 492854
rect 527866 492618 528102 492854
rect 527546 456938 527782 457174
rect 527866 456938 528102 457174
rect 527546 456618 527782 456854
rect 527866 456618 528102 456854
rect 527546 420938 527782 421174
rect 527866 420938 528102 421174
rect 527546 420618 527782 420854
rect 527866 420618 528102 420854
rect 527546 384938 527782 385174
rect 527866 384938 528102 385174
rect 527546 384618 527782 384854
rect 527866 384618 528102 384854
rect 527546 348938 527782 349174
rect 527866 348938 528102 349174
rect 527546 348618 527782 348854
rect 527866 348618 528102 348854
rect 527546 312938 527782 313174
rect 527866 312938 528102 313174
rect 527546 312618 527782 312854
rect 527866 312618 528102 312854
rect 527546 276938 527782 277174
rect 527866 276938 528102 277174
rect 527546 276618 527782 276854
rect 527866 276618 528102 276854
rect 527546 240938 527782 241174
rect 527866 240938 528102 241174
rect 527546 240618 527782 240854
rect 527866 240618 528102 240854
rect 527546 204938 527782 205174
rect 527866 204938 528102 205174
rect 527546 204618 527782 204854
rect 527866 204618 528102 204854
rect 527546 168938 527782 169174
rect 527866 168938 528102 169174
rect 527546 168618 527782 168854
rect 527866 168618 528102 168854
rect 527546 132938 527782 133174
rect 527866 132938 528102 133174
rect 527546 132618 527782 132854
rect 527866 132618 528102 132854
rect 527546 96938 527782 97174
rect 527866 96938 528102 97174
rect 527546 96618 527782 96854
rect 527866 96618 528102 96854
rect 527546 60938 527782 61174
rect 527866 60938 528102 61174
rect 527546 60618 527782 60854
rect 527866 60618 528102 60854
rect 527546 24938 527782 25174
rect 527866 24938 528102 25174
rect 527546 24618 527782 24854
rect 527866 24618 528102 24854
rect 527546 -3462 527782 -3226
rect 527866 -3462 528102 -3226
rect 527546 -3782 527782 -3546
rect 527866 -3782 528102 -3546
rect 531266 676658 531502 676894
rect 531586 676658 531822 676894
rect 531266 676338 531502 676574
rect 531586 676338 531822 676574
rect 531266 640658 531502 640894
rect 531586 640658 531822 640894
rect 531266 640338 531502 640574
rect 531586 640338 531822 640574
rect 531266 604658 531502 604894
rect 531586 604658 531822 604894
rect 531266 604338 531502 604574
rect 531586 604338 531822 604574
rect 531266 568658 531502 568894
rect 531586 568658 531822 568894
rect 531266 568338 531502 568574
rect 531586 568338 531822 568574
rect 531266 532658 531502 532894
rect 531586 532658 531822 532894
rect 531266 532338 531502 532574
rect 531586 532338 531822 532574
rect 531266 496658 531502 496894
rect 531586 496658 531822 496894
rect 531266 496338 531502 496574
rect 531586 496338 531822 496574
rect 531266 460658 531502 460894
rect 531586 460658 531822 460894
rect 531266 460338 531502 460574
rect 531586 460338 531822 460574
rect 531266 424658 531502 424894
rect 531586 424658 531822 424894
rect 531266 424338 531502 424574
rect 531586 424338 531822 424574
rect 531266 388658 531502 388894
rect 531586 388658 531822 388894
rect 531266 388338 531502 388574
rect 531586 388338 531822 388574
rect 531266 352658 531502 352894
rect 531586 352658 531822 352894
rect 531266 352338 531502 352574
rect 531586 352338 531822 352574
rect 531266 316658 531502 316894
rect 531586 316658 531822 316894
rect 531266 316338 531502 316574
rect 531586 316338 531822 316574
rect 531266 280658 531502 280894
rect 531586 280658 531822 280894
rect 531266 280338 531502 280574
rect 531586 280338 531822 280574
rect 531266 244658 531502 244894
rect 531586 244658 531822 244894
rect 531266 244338 531502 244574
rect 531586 244338 531822 244574
rect 531266 208658 531502 208894
rect 531586 208658 531822 208894
rect 531266 208338 531502 208574
rect 531586 208338 531822 208574
rect 531266 172658 531502 172894
rect 531586 172658 531822 172894
rect 531266 172338 531502 172574
rect 531586 172338 531822 172574
rect 531266 136658 531502 136894
rect 531586 136658 531822 136894
rect 531266 136338 531502 136574
rect 531586 136338 531822 136574
rect 531266 100658 531502 100894
rect 531586 100658 531822 100894
rect 531266 100338 531502 100574
rect 531586 100338 531822 100574
rect 531266 64658 531502 64894
rect 531586 64658 531822 64894
rect 531266 64338 531502 64574
rect 531586 64338 531822 64574
rect 531266 28658 531502 28894
rect 531586 28658 531822 28894
rect 531266 28338 531502 28574
rect 531586 28338 531822 28574
rect 531266 -5382 531502 -5146
rect 531586 -5382 531822 -5146
rect 531266 -5702 531502 -5466
rect 531586 -5702 531822 -5466
rect 552986 710362 553222 710598
rect 553306 710362 553542 710598
rect 552986 710042 553222 710278
rect 553306 710042 553542 710278
rect 549266 708442 549502 708678
rect 549586 708442 549822 708678
rect 549266 708122 549502 708358
rect 549586 708122 549822 708358
rect 545546 706522 545782 706758
rect 545866 706522 546102 706758
rect 545546 706202 545782 706438
rect 545866 706202 546102 706438
rect 534986 680378 535222 680614
rect 535306 680378 535542 680614
rect 534986 680058 535222 680294
rect 535306 680058 535542 680294
rect 534986 644378 535222 644614
rect 535306 644378 535542 644614
rect 534986 644058 535222 644294
rect 535306 644058 535542 644294
rect 534986 608378 535222 608614
rect 535306 608378 535542 608614
rect 534986 608058 535222 608294
rect 535306 608058 535542 608294
rect 534986 572378 535222 572614
rect 535306 572378 535542 572614
rect 534986 572058 535222 572294
rect 535306 572058 535542 572294
rect 534986 536378 535222 536614
rect 535306 536378 535542 536614
rect 534986 536058 535222 536294
rect 535306 536058 535542 536294
rect 534986 500378 535222 500614
rect 535306 500378 535542 500614
rect 534986 500058 535222 500294
rect 535306 500058 535542 500294
rect 534986 464378 535222 464614
rect 535306 464378 535542 464614
rect 534986 464058 535222 464294
rect 535306 464058 535542 464294
rect 534986 428378 535222 428614
rect 535306 428378 535542 428614
rect 534986 428058 535222 428294
rect 535306 428058 535542 428294
rect 534986 392378 535222 392614
rect 535306 392378 535542 392614
rect 534986 392058 535222 392294
rect 535306 392058 535542 392294
rect 534986 356378 535222 356614
rect 535306 356378 535542 356614
rect 534986 356058 535222 356294
rect 535306 356058 535542 356294
rect 534986 320378 535222 320614
rect 535306 320378 535542 320614
rect 534986 320058 535222 320294
rect 535306 320058 535542 320294
rect 534986 284378 535222 284614
rect 535306 284378 535542 284614
rect 534986 284058 535222 284294
rect 535306 284058 535542 284294
rect 534986 248378 535222 248614
rect 535306 248378 535542 248614
rect 534986 248058 535222 248294
rect 535306 248058 535542 248294
rect 534986 212378 535222 212614
rect 535306 212378 535542 212614
rect 534986 212058 535222 212294
rect 535306 212058 535542 212294
rect 534986 176378 535222 176614
rect 535306 176378 535542 176614
rect 534986 176058 535222 176294
rect 535306 176058 535542 176294
rect 534986 140378 535222 140614
rect 535306 140378 535542 140614
rect 534986 140058 535222 140294
rect 535306 140058 535542 140294
rect 534986 104378 535222 104614
rect 535306 104378 535542 104614
rect 534986 104058 535222 104294
rect 535306 104058 535542 104294
rect 534986 68378 535222 68614
rect 535306 68378 535542 68614
rect 534986 68058 535222 68294
rect 535306 68058 535542 68294
rect 534986 32378 535222 32614
rect 535306 32378 535542 32614
rect 534986 32058 535222 32294
rect 535306 32058 535542 32294
rect 516986 -6342 517222 -6106
rect 517306 -6342 517542 -6106
rect 516986 -6662 517222 -6426
rect 517306 -6662 517542 -6426
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 690938 545782 691174
rect 545866 690938 546102 691174
rect 545546 690618 545782 690854
rect 545866 690618 546102 690854
rect 545546 654938 545782 655174
rect 545866 654938 546102 655174
rect 545546 654618 545782 654854
rect 545866 654618 546102 654854
rect 545546 618938 545782 619174
rect 545866 618938 546102 619174
rect 545546 618618 545782 618854
rect 545866 618618 546102 618854
rect 545546 582938 545782 583174
rect 545866 582938 546102 583174
rect 545546 582618 545782 582854
rect 545866 582618 546102 582854
rect 545546 546938 545782 547174
rect 545866 546938 546102 547174
rect 545546 546618 545782 546854
rect 545866 546618 546102 546854
rect 545546 510938 545782 511174
rect 545866 510938 546102 511174
rect 545546 510618 545782 510854
rect 545866 510618 546102 510854
rect 545546 474938 545782 475174
rect 545866 474938 546102 475174
rect 545546 474618 545782 474854
rect 545866 474618 546102 474854
rect 545546 438938 545782 439174
rect 545866 438938 546102 439174
rect 545546 438618 545782 438854
rect 545866 438618 546102 438854
rect 545546 402938 545782 403174
rect 545866 402938 546102 403174
rect 545546 402618 545782 402854
rect 545866 402618 546102 402854
rect 545546 366938 545782 367174
rect 545866 366938 546102 367174
rect 545546 366618 545782 366854
rect 545866 366618 546102 366854
rect 545546 330938 545782 331174
rect 545866 330938 546102 331174
rect 545546 330618 545782 330854
rect 545866 330618 546102 330854
rect 545546 294938 545782 295174
rect 545866 294938 546102 295174
rect 545546 294618 545782 294854
rect 545866 294618 546102 294854
rect 545546 258938 545782 259174
rect 545866 258938 546102 259174
rect 545546 258618 545782 258854
rect 545866 258618 546102 258854
rect 545546 222938 545782 223174
rect 545866 222938 546102 223174
rect 545546 222618 545782 222854
rect 545866 222618 546102 222854
rect 545546 186938 545782 187174
rect 545866 186938 546102 187174
rect 545546 186618 545782 186854
rect 545866 186618 546102 186854
rect 545546 150938 545782 151174
rect 545866 150938 546102 151174
rect 545546 150618 545782 150854
rect 545866 150618 546102 150854
rect 545546 114938 545782 115174
rect 545866 114938 546102 115174
rect 545546 114618 545782 114854
rect 545866 114618 546102 114854
rect 545546 78938 545782 79174
rect 545866 78938 546102 79174
rect 545546 78618 545782 78854
rect 545866 78618 546102 78854
rect 545546 42938 545782 43174
rect 545866 42938 546102 43174
rect 545546 42618 545782 42854
rect 545866 42618 546102 42854
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -2502 545782 -2266
rect 545866 -2502 546102 -2266
rect 545546 -2822 545782 -2586
rect 545866 -2822 546102 -2586
rect 549266 694658 549502 694894
rect 549586 694658 549822 694894
rect 549266 694338 549502 694574
rect 549586 694338 549822 694574
rect 549266 658658 549502 658894
rect 549586 658658 549822 658894
rect 549266 658338 549502 658574
rect 549586 658338 549822 658574
rect 549266 622658 549502 622894
rect 549586 622658 549822 622894
rect 549266 622338 549502 622574
rect 549586 622338 549822 622574
rect 549266 586658 549502 586894
rect 549586 586658 549822 586894
rect 549266 586338 549502 586574
rect 549586 586338 549822 586574
rect 549266 550658 549502 550894
rect 549586 550658 549822 550894
rect 549266 550338 549502 550574
rect 549586 550338 549822 550574
rect 549266 514658 549502 514894
rect 549586 514658 549822 514894
rect 549266 514338 549502 514574
rect 549586 514338 549822 514574
rect 549266 478658 549502 478894
rect 549586 478658 549822 478894
rect 549266 478338 549502 478574
rect 549586 478338 549822 478574
rect 549266 442658 549502 442894
rect 549586 442658 549822 442894
rect 549266 442338 549502 442574
rect 549586 442338 549822 442574
rect 549266 406658 549502 406894
rect 549586 406658 549822 406894
rect 549266 406338 549502 406574
rect 549586 406338 549822 406574
rect 549266 370658 549502 370894
rect 549586 370658 549822 370894
rect 549266 370338 549502 370574
rect 549586 370338 549822 370574
rect 549266 334658 549502 334894
rect 549586 334658 549822 334894
rect 549266 334338 549502 334574
rect 549586 334338 549822 334574
rect 549266 298658 549502 298894
rect 549586 298658 549822 298894
rect 549266 298338 549502 298574
rect 549586 298338 549822 298574
rect 549266 262658 549502 262894
rect 549586 262658 549822 262894
rect 549266 262338 549502 262574
rect 549586 262338 549822 262574
rect 549266 226658 549502 226894
rect 549586 226658 549822 226894
rect 549266 226338 549502 226574
rect 549586 226338 549822 226574
rect 549266 190658 549502 190894
rect 549586 190658 549822 190894
rect 549266 190338 549502 190574
rect 549586 190338 549822 190574
rect 549266 154658 549502 154894
rect 549586 154658 549822 154894
rect 549266 154338 549502 154574
rect 549586 154338 549822 154574
rect 549266 118658 549502 118894
rect 549586 118658 549822 118894
rect 549266 118338 549502 118574
rect 549586 118338 549822 118574
rect 549266 82658 549502 82894
rect 549586 82658 549822 82894
rect 549266 82338 549502 82574
rect 549586 82338 549822 82574
rect 549266 46658 549502 46894
rect 549586 46658 549822 46894
rect 549266 46338 549502 46574
rect 549586 46338 549822 46574
rect 549266 10658 549502 10894
rect 549586 10658 549822 10894
rect 549266 10338 549502 10574
rect 549586 10338 549822 10574
rect 549266 -4422 549502 -4186
rect 549586 -4422 549822 -4186
rect 549266 -4742 549502 -4506
rect 549586 -4742 549822 -4506
rect 570986 711322 571222 711558
rect 571306 711322 571542 711558
rect 570986 711002 571222 711238
rect 571306 711002 571542 711238
rect 567266 709402 567502 709638
rect 567586 709402 567822 709638
rect 567266 709082 567502 709318
rect 567586 709082 567822 709318
rect 563546 707482 563782 707718
rect 563866 707482 564102 707718
rect 563546 707162 563782 707398
rect 563866 707162 564102 707398
rect 552986 698378 553222 698614
rect 553306 698378 553542 698614
rect 552986 698058 553222 698294
rect 553306 698058 553542 698294
rect 552986 662378 553222 662614
rect 553306 662378 553542 662614
rect 552986 662058 553222 662294
rect 553306 662058 553542 662294
rect 552986 626378 553222 626614
rect 553306 626378 553542 626614
rect 552986 626058 553222 626294
rect 553306 626058 553542 626294
rect 552986 590378 553222 590614
rect 553306 590378 553542 590614
rect 552986 590058 553222 590294
rect 553306 590058 553542 590294
rect 552986 554378 553222 554614
rect 553306 554378 553542 554614
rect 552986 554058 553222 554294
rect 553306 554058 553542 554294
rect 552986 518378 553222 518614
rect 553306 518378 553542 518614
rect 552986 518058 553222 518294
rect 553306 518058 553542 518294
rect 552986 482378 553222 482614
rect 553306 482378 553542 482614
rect 552986 482058 553222 482294
rect 553306 482058 553542 482294
rect 552986 446378 553222 446614
rect 553306 446378 553542 446614
rect 552986 446058 553222 446294
rect 553306 446058 553542 446294
rect 552986 410378 553222 410614
rect 553306 410378 553542 410614
rect 552986 410058 553222 410294
rect 553306 410058 553542 410294
rect 552986 374378 553222 374614
rect 553306 374378 553542 374614
rect 552986 374058 553222 374294
rect 553306 374058 553542 374294
rect 552986 338378 553222 338614
rect 553306 338378 553542 338614
rect 552986 338058 553222 338294
rect 553306 338058 553542 338294
rect 552986 302378 553222 302614
rect 553306 302378 553542 302614
rect 552986 302058 553222 302294
rect 553306 302058 553542 302294
rect 552986 266378 553222 266614
rect 553306 266378 553542 266614
rect 552986 266058 553222 266294
rect 553306 266058 553542 266294
rect 552986 230378 553222 230614
rect 553306 230378 553542 230614
rect 552986 230058 553222 230294
rect 553306 230058 553542 230294
rect 552986 194378 553222 194614
rect 553306 194378 553542 194614
rect 552986 194058 553222 194294
rect 553306 194058 553542 194294
rect 552986 158378 553222 158614
rect 553306 158378 553542 158614
rect 552986 158058 553222 158294
rect 553306 158058 553542 158294
rect 552986 122378 553222 122614
rect 553306 122378 553542 122614
rect 552986 122058 553222 122294
rect 553306 122058 553542 122294
rect 552986 86378 553222 86614
rect 553306 86378 553542 86614
rect 552986 86058 553222 86294
rect 553306 86058 553542 86294
rect 552986 50378 553222 50614
rect 553306 50378 553542 50614
rect 552986 50058 553222 50294
rect 553306 50058 553542 50294
rect 552986 14378 553222 14614
rect 553306 14378 553542 14614
rect 552986 14058 553222 14294
rect 553306 14058 553542 14294
rect 534986 -7302 535222 -7066
rect 535306 -7302 535542 -7066
rect 534986 -7622 535222 -7386
rect 535306 -7622 535542 -7386
rect 559826 705562 560062 705798
rect 560146 705562 560382 705798
rect 559826 705242 560062 705478
rect 560146 705242 560382 705478
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -1542 560062 -1306
rect 560146 -1542 560382 -1306
rect 559826 -1862 560062 -1626
rect 560146 -1862 560382 -1626
rect 563546 672938 563782 673174
rect 563866 672938 564102 673174
rect 563546 672618 563782 672854
rect 563866 672618 564102 672854
rect 563546 636938 563782 637174
rect 563866 636938 564102 637174
rect 563546 636618 563782 636854
rect 563866 636618 564102 636854
rect 563546 600938 563782 601174
rect 563866 600938 564102 601174
rect 563546 600618 563782 600854
rect 563866 600618 564102 600854
rect 563546 564938 563782 565174
rect 563866 564938 564102 565174
rect 563546 564618 563782 564854
rect 563866 564618 564102 564854
rect 563546 528938 563782 529174
rect 563866 528938 564102 529174
rect 563546 528618 563782 528854
rect 563866 528618 564102 528854
rect 563546 492938 563782 493174
rect 563866 492938 564102 493174
rect 563546 492618 563782 492854
rect 563866 492618 564102 492854
rect 563546 456938 563782 457174
rect 563866 456938 564102 457174
rect 563546 456618 563782 456854
rect 563866 456618 564102 456854
rect 563546 420938 563782 421174
rect 563866 420938 564102 421174
rect 563546 420618 563782 420854
rect 563866 420618 564102 420854
rect 563546 384938 563782 385174
rect 563866 384938 564102 385174
rect 563546 384618 563782 384854
rect 563866 384618 564102 384854
rect 563546 348938 563782 349174
rect 563866 348938 564102 349174
rect 563546 348618 563782 348854
rect 563866 348618 564102 348854
rect 563546 312938 563782 313174
rect 563866 312938 564102 313174
rect 563546 312618 563782 312854
rect 563866 312618 564102 312854
rect 563546 276938 563782 277174
rect 563866 276938 564102 277174
rect 563546 276618 563782 276854
rect 563866 276618 564102 276854
rect 563546 240938 563782 241174
rect 563866 240938 564102 241174
rect 563546 240618 563782 240854
rect 563866 240618 564102 240854
rect 563546 204938 563782 205174
rect 563866 204938 564102 205174
rect 563546 204618 563782 204854
rect 563866 204618 564102 204854
rect 563546 168938 563782 169174
rect 563866 168938 564102 169174
rect 563546 168618 563782 168854
rect 563866 168618 564102 168854
rect 563546 132938 563782 133174
rect 563866 132938 564102 133174
rect 563546 132618 563782 132854
rect 563866 132618 564102 132854
rect 563546 96938 563782 97174
rect 563866 96938 564102 97174
rect 563546 96618 563782 96854
rect 563866 96618 564102 96854
rect 563546 60938 563782 61174
rect 563866 60938 564102 61174
rect 563546 60618 563782 60854
rect 563866 60618 564102 60854
rect 563546 24938 563782 25174
rect 563866 24938 564102 25174
rect 563546 24618 563782 24854
rect 563866 24618 564102 24854
rect 563546 -3462 563782 -3226
rect 563866 -3462 564102 -3226
rect 563546 -3782 563782 -3546
rect 563866 -3782 564102 -3546
rect 567266 676658 567502 676894
rect 567586 676658 567822 676894
rect 567266 676338 567502 676574
rect 567586 676338 567822 676574
rect 567266 640658 567502 640894
rect 567586 640658 567822 640894
rect 567266 640338 567502 640574
rect 567586 640338 567822 640574
rect 567266 604658 567502 604894
rect 567586 604658 567822 604894
rect 567266 604338 567502 604574
rect 567586 604338 567822 604574
rect 567266 568658 567502 568894
rect 567586 568658 567822 568894
rect 567266 568338 567502 568574
rect 567586 568338 567822 568574
rect 567266 532658 567502 532894
rect 567586 532658 567822 532894
rect 567266 532338 567502 532574
rect 567586 532338 567822 532574
rect 567266 496658 567502 496894
rect 567586 496658 567822 496894
rect 567266 496338 567502 496574
rect 567586 496338 567822 496574
rect 567266 460658 567502 460894
rect 567586 460658 567822 460894
rect 567266 460338 567502 460574
rect 567586 460338 567822 460574
rect 567266 424658 567502 424894
rect 567586 424658 567822 424894
rect 567266 424338 567502 424574
rect 567586 424338 567822 424574
rect 567266 388658 567502 388894
rect 567586 388658 567822 388894
rect 567266 388338 567502 388574
rect 567586 388338 567822 388574
rect 567266 352658 567502 352894
rect 567586 352658 567822 352894
rect 567266 352338 567502 352574
rect 567586 352338 567822 352574
rect 567266 316658 567502 316894
rect 567586 316658 567822 316894
rect 567266 316338 567502 316574
rect 567586 316338 567822 316574
rect 567266 280658 567502 280894
rect 567586 280658 567822 280894
rect 567266 280338 567502 280574
rect 567586 280338 567822 280574
rect 567266 244658 567502 244894
rect 567586 244658 567822 244894
rect 567266 244338 567502 244574
rect 567586 244338 567822 244574
rect 567266 208658 567502 208894
rect 567586 208658 567822 208894
rect 567266 208338 567502 208574
rect 567586 208338 567822 208574
rect 567266 172658 567502 172894
rect 567586 172658 567822 172894
rect 567266 172338 567502 172574
rect 567586 172338 567822 172574
rect 567266 136658 567502 136894
rect 567586 136658 567822 136894
rect 567266 136338 567502 136574
rect 567586 136338 567822 136574
rect 567266 100658 567502 100894
rect 567586 100658 567822 100894
rect 567266 100338 567502 100574
rect 567586 100338 567822 100574
rect 567266 64658 567502 64894
rect 567586 64658 567822 64894
rect 567266 64338 567502 64574
rect 567586 64338 567822 64574
rect 567266 28658 567502 28894
rect 567586 28658 567822 28894
rect 567266 28338 567502 28574
rect 567586 28338 567822 28574
rect 567266 -5382 567502 -5146
rect 567586 -5382 567822 -5146
rect 567266 -5702 567502 -5466
rect 567586 -5702 567822 -5466
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 581546 706522 581782 706758
rect 581866 706522 582102 706758
rect 581546 706202 581782 706438
rect 581866 706202 582102 706438
rect 570986 680378 571222 680614
rect 571306 680378 571542 680614
rect 570986 680058 571222 680294
rect 571306 680058 571542 680294
rect 570986 644378 571222 644614
rect 571306 644378 571542 644614
rect 570986 644058 571222 644294
rect 571306 644058 571542 644294
rect 570986 608378 571222 608614
rect 571306 608378 571542 608614
rect 570986 608058 571222 608294
rect 571306 608058 571542 608294
rect 570986 572378 571222 572614
rect 571306 572378 571542 572614
rect 570986 572058 571222 572294
rect 571306 572058 571542 572294
rect 570986 536378 571222 536614
rect 571306 536378 571542 536614
rect 570986 536058 571222 536294
rect 571306 536058 571542 536294
rect 570986 500378 571222 500614
rect 571306 500378 571542 500614
rect 570986 500058 571222 500294
rect 571306 500058 571542 500294
rect 570986 464378 571222 464614
rect 571306 464378 571542 464614
rect 570986 464058 571222 464294
rect 571306 464058 571542 464294
rect 570986 428378 571222 428614
rect 571306 428378 571542 428614
rect 570986 428058 571222 428294
rect 571306 428058 571542 428294
rect 570986 392378 571222 392614
rect 571306 392378 571542 392614
rect 570986 392058 571222 392294
rect 571306 392058 571542 392294
rect 570986 356378 571222 356614
rect 571306 356378 571542 356614
rect 570986 356058 571222 356294
rect 571306 356058 571542 356294
rect 570986 320378 571222 320614
rect 571306 320378 571542 320614
rect 570986 320058 571222 320294
rect 571306 320058 571542 320294
rect 570986 284378 571222 284614
rect 571306 284378 571542 284614
rect 570986 284058 571222 284294
rect 571306 284058 571542 284294
rect 570986 248378 571222 248614
rect 571306 248378 571542 248614
rect 570986 248058 571222 248294
rect 571306 248058 571542 248294
rect 570986 212378 571222 212614
rect 571306 212378 571542 212614
rect 570986 212058 571222 212294
rect 571306 212058 571542 212294
rect 570986 176378 571222 176614
rect 571306 176378 571542 176614
rect 570986 176058 571222 176294
rect 571306 176058 571542 176294
rect 570986 140378 571222 140614
rect 571306 140378 571542 140614
rect 570986 140058 571222 140294
rect 571306 140058 571542 140294
rect 570986 104378 571222 104614
rect 571306 104378 571542 104614
rect 570986 104058 571222 104294
rect 571306 104058 571542 104294
rect 570986 68378 571222 68614
rect 571306 68378 571542 68614
rect 570986 68058 571222 68294
rect 571306 68058 571542 68294
rect 570986 32378 571222 32614
rect 571306 32378 571542 32614
rect 570986 32058 571222 32294
rect 571306 32058 571542 32294
rect 552986 -6342 553222 -6106
rect 553306 -6342 553542 -6106
rect 552986 -6662 553222 -6426
rect 553306 -6662 553542 -6426
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 669218 586538 669454
rect 586622 669218 586858 669454
rect 586302 668898 586538 669134
rect 586622 668898 586858 669134
rect 586302 633218 586538 633454
rect 586622 633218 586858 633454
rect 586302 632898 586538 633134
rect 586622 632898 586858 633134
rect 586302 597218 586538 597454
rect 586622 597218 586858 597454
rect 586302 596898 586538 597134
rect 586622 596898 586858 597134
rect 586302 561218 586538 561454
rect 586622 561218 586858 561454
rect 586302 560898 586538 561134
rect 586622 560898 586858 561134
rect 586302 525218 586538 525454
rect 586622 525218 586858 525454
rect 586302 524898 586538 525134
rect 586622 524898 586858 525134
rect 586302 489218 586538 489454
rect 586622 489218 586858 489454
rect 586302 488898 586538 489134
rect 586622 488898 586858 489134
rect 586302 453218 586538 453454
rect 586622 453218 586858 453454
rect 586302 452898 586538 453134
rect 586622 452898 586858 453134
rect 586302 417218 586538 417454
rect 586622 417218 586858 417454
rect 586302 416898 586538 417134
rect 586622 416898 586858 417134
rect 586302 381218 586538 381454
rect 586622 381218 586858 381454
rect 586302 380898 586538 381134
rect 586622 380898 586858 381134
rect 586302 345218 586538 345454
rect 586622 345218 586858 345454
rect 586302 344898 586538 345134
rect 586622 344898 586858 345134
rect 586302 309218 586538 309454
rect 586622 309218 586858 309454
rect 586302 308898 586538 309134
rect 586622 308898 586858 309134
rect 586302 273218 586538 273454
rect 586622 273218 586858 273454
rect 586302 272898 586538 273134
rect 586622 272898 586858 273134
rect 586302 237218 586538 237454
rect 586622 237218 586858 237454
rect 586302 236898 586538 237134
rect 586622 236898 586858 237134
rect 586302 201218 586538 201454
rect 586622 201218 586858 201454
rect 586302 200898 586538 201134
rect 586622 200898 586858 201134
rect 586302 165218 586538 165454
rect 586622 165218 586858 165454
rect 586302 164898 586538 165134
rect 586622 164898 586858 165134
rect 586302 129218 586538 129454
rect 586622 129218 586858 129454
rect 586302 128898 586538 129134
rect 586622 128898 586858 129134
rect 586302 93218 586538 93454
rect 586622 93218 586858 93454
rect 586302 92898 586538 93134
rect 586622 92898 586858 93134
rect 586302 57218 586538 57454
rect 586622 57218 586858 57454
rect 586302 56898 586538 57134
rect 586622 56898 586858 57134
rect 586302 21218 586538 21454
rect 586622 21218 586858 21454
rect 586302 20898 586538 21134
rect 586622 20898 586858 21134
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 690938 587498 691174
rect 587582 690938 587818 691174
rect 587262 690618 587498 690854
rect 587582 690618 587818 690854
rect 587262 654938 587498 655174
rect 587582 654938 587818 655174
rect 587262 654618 587498 654854
rect 587582 654618 587818 654854
rect 587262 618938 587498 619174
rect 587582 618938 587818 619174
rect 587262 618618 587498 618854
rect 587582 618618 587818 618854
rect 587262 582938 587498 583174
rect 587582 582938 587818 583174
rect 587262 582618 587498 582854
rect 587582 582618 587818 582854
rect 587262 546938 587498 547174
rect 587582 546938 587818 547174
rect 587262 546618 587498 546854
rect 587582 546618 587818 546854
rect 587262 510938 587498 511174
rect 587582 510938 587818 511174
rect 587262 510618 587498 510854
rect 587582 510618 587818 510854
rect 587262 474938 587498 475174
rect 587582 474938 587818 475174
rect 587262 474618 587498 474854
rect 587582 474618 587818 474854
rect 587262 438938 587498 439174
rect 587582 438938 587818 439174
rect 587262 438618 587498 438854
rect 587582 438618 587818 438854
rect 587262 402938 587498 403174
rect 587582 402938 587818 403174
rect 587262 402618 587498 402854
rect 587582 402618 587818 402854
rect 587262 366938 587498 367174
rect 587582 366938 587818 367174
rect 587262 366618 587498 366854
rect 587582 366618 587818 366854
rect 587262 330938 587498 331174
rect 587582 330938 587818 331174
rect 587262 330618 587498 330854
rect 587582 330618 587818 330854
rect 587262 294938 587498 295174
rect 587582 294938 587818 295174
rect 587262 294618 587498 294854
rect 587582 294618 587818 294854
rect 587262 258938 587498 259174
rect 587582 258938 587818 259174
rect 587262 258618 587498 258854
rect 587582 258618 587818 258854
rect 587262 222938 587498 223174
rect 587582 222938 587818 223174
rect 587262 222618 587498 222854
rect 587582 222618 587818 222854
rect 587262 186938 587498 187174
rect 587582 186938 587818 187174
rect 587262 186618 587498 186854
rect 587582 186618 587818 186854
rect 587262 150938 587498 151174
rect 587582 150938 587818 151174
rect 587262 150618 587498 150854
rect 587582 150618 587818 150854
rect 587262 114938 587498 115174
rect 587582 114938 587818 115174
rect 587262 114618 587498 114854
rect 587582 114618 587818 114854
rect 587262 78938 587498 79174
rect 587582 78938 587818 79174
rect 587262 78618 587498 78854
rect 587582 78618 587818 78854
rect 587262 42938 587498 43174
rect 587582 42938 587818 43174
rect 587262 42618 587498 42854
rect 587582 42618 587818 42854
rect 587262 6938 587498 7174
rect 587582 6938 587818 7174
rect 587262 6618 587498 6854
rect 587582 6618 587818 6854
rect 581546 -2502 581782 -2266
rect 581866 -2502 582102 -2266
rect 581546 -2822 581782 -2586
rect 581866 -2822 582102 -2586
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 672938 588458 673174
rect 588542 672938 588778 673174
rect 588222 672618 588458 672854
rect 588542 672618 588778 672854
rect 588222 636938 588458 637174
rect 588542 636938 588778 637174
rect 588222 636618 588458 636854
rect 588542 636618 588778 636854
rect 588222 600938 588458 601174
rect 588542 600938 588778 601174
rect 588222 600618 588458 600854
rect 588542 600618 588778 600854
rect 588222 564938 588458 565174
rect 588542 564938 588778 565174
rect 588222 564618 588458 564854
rect 588542 564618 588778 564854
rect 588222 528938 588458 529174
rect 588542 528938 588778 529174
rect 588222 528618 588458 528854
rect 588542 528618 588778 528854
rect 588222 492938 588458 493174
rect 588542 492938 588778 493174
rect 588222 492618 588458 492854
rect 588542 492618 588778 492854
rect 588222 456938 588458 457174
rect 588542 456938 588778 457174
rect 588222 456618 588458 456854
rect 588542 456618 588778 456854
rect 588222 420938 588458 421174
rect 588542 420938 588778 421174
rect 588222 420618 588458 420854
rect 588542 420618 588778 420854
rect 588222 384938 588458 385174
rect 588542 384938 588778 385174
rect 588222 384618 588458 384854
rect 588542 384618 588778 384854
rect 588222 348938 588458 349174
rect 588542 348938 588778 349174
rect 588222 348618 588458 348854
rect 588542 348618 588778 348854
rect 588222 312938 588458 313174
rect 588542 312938 588778 313174
rect 588222 312618 588458 312854
rect 588542 312618 588778 312854
rect 588222 276938 588458 277174
rect 588542 276938 588778 277174
rect 588222 276618 588458 276854
rect 588542 276618 588778 276854
rect 588222 240938 588458 241174
rect 588542 240938 588778 241174
rect 588222 240618 588458 240854
rect 588542 240618 588778 240854
rect 588222 204938 588458 205174
rect 588542 204938 588778 205174
rect 588222 204618 588458 204854
rect 588542 204618 588778 204854
rect 588222 168938 588458 169174
rect 588542 168938 588778 169174
rect 588222 168618 588458 168854
rect 588542 168618 588778 168854
rect 588222 132938 588458 133174
rect 588542 132938 588778 133174
rect 588222 132618 588458 132854
rect 588542 132618 588778 132854
rect 588222 96938 588458 97174
rect 588542 96938 588778 97174
rect 588222 96618 588458 96854
rect 588542 96618 588778 96854
rect 588222 60938 588458 61174
rect 588542 60938 588778 61174
rect 588222 60618 588458 60854
rect 588542 60618 588778 60854
rect 588222 24938 588458 25174
rect 588542 24938 588778 25174
rect 588222 24618 588458 24854
rect 588542 24618 588778 24854
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 694658 589418 694894
rect 589502 694658 589738 694894
rect 589182 694338 589418 694574
rect 589502 694338 589738 694574
rect 589182 658658 589418 658894
rect 589502 658658 589738 658894
rect 589182 658338 589418 658574
rect 589502 658338 589738 658574
rect 589182 622658 589418 622894
rect 589502 622658 589738 622894
rect 589182 622338 589418 622574
rect 589502 622338 589738 622574
rect 589182 586658 589418 586894
rect 589502 586658 589738 586894
rect 589182 586338 589418 586574
rect 589502 586338 589738 586574
rect 589182 550658 589418 550894
rect 589502 550658 589738 550894
rect 589182 550338 589418 550574
rect 589502 550338 589738 550574
rect 589182 514658 589418 514894
rect 589502 514658 589738 514894
rect 589182 514338 589418 514574
rect 589502 514338 589738 514574
rect 589182 478658 589418 478894
rect 589502 478658 589738 478894
rect 589182 478338 589418 478574
rect 589502 478338 589738 478574
rect 589182 442658 589418 442894
rect 589502 442658 589738 442894
rect 589182 442338 589418 442574
rect 589502 442338 589738 442574
rect 589182 406658 589418 406894
rect 589502 406658 589738 406894
rect 589182 406338 589418 406574
rect 589502 406338 589738 406574
rect 589182 370658 589418 370894
rect 589502 370658 589738 370894
rect 589182 370338 589418 370574
rect 589502 370338 589738 370574
rect 589182 334658 589418 334894
rect 589502 334658 589738 334894
rect 589182 334338 589418 334574
rect 589502 334338 589738 334574
rect 589182 298658 589418 298894
rect 589502 298658 589738 298894
rect 589182 298338 589418 298574
rect 589502 298338 589738 298574
rect 589182 262658 589418 262894
rect 589502 262658 589738 262894
rect 589182 262338 589418 262574
rect 589502 262338 589738 262574
rect 589182 226658 589418 226894
rect 589502 226658 589738 226894
rect 589182 226338 589418 226574
rect 589502 226338 589738 226574
rect 589182 190658 589418 190894
rect 589502 190658 589738 190894
rect 589182 190338 589418 190574
rect 589502 190338 589738 190574
rect 589182 154658 589418 154894
rect 589502 154658 589738 154894
rect 589182 154338 589418 154574
rect 589502 154338 589738 154574
rect 589182 118658 589418 118894
rect 589502 118658 589738 118894
rect 589182 118338 589418 118574
rect 589502 118338 589738 118574
rect 589182 82658 589418 82894
rect 589502 82658 589738 82894
rect 589182 82338 589418 82574
rect 589502 82338 589738 82574
rect 589182 46658 589418 46894
rect 589502 46658 589738 46894
rect 589182 46338 589418 46574
rect 589502 46338 589738 46574
rect 589182 10658 589418 10894
rect 589502 10658 589738 10894
rect 589182 10338 589418 10574
rect 589502 10338 589738 10574
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 676658 590378 676894
rect 590462 676658 590698 676894
rect 590142 676338 590378 676574
rect 590462 676338 590698 676574
rect 590142 640658 590378 640894
rect 590462 640658 590698 640894
rect 590142 640338 590378 640574
rect 590462 640338 590698 640574
rect 590142 604658 590378 604894
rect 590462 604658 590698 604894
rect 590142 604338 590378 604574
rect 590462 604338 590698 604574
rect 590142 568658 590378 568894
rect 590462 568658 590698 568894
rect 590142 568338 590378 568574
rect 590462 568338 590698 568574
rect 590142 532658 590378 532894
rect 590462 532658 590698 532894
rect 590142 532338 590378 532574
rect 590462 532338 590698 532574
rect 590142 496658 590378 496894
rect 590462 496658 590698 496894
rect 590142 496338 590378 496574
rect 590462 496338 590698 496574
rect 590142 460658 590378 460894
rect 590462 460658 590698 460894
rect 590142 460338 590378 460574
rect 590462 460338 590698 460574
rect 590142 424658 590378 424894
rect 590462 424658 590698 424894
rect 590142 424338 590378 424574
rect 590462 424338 590698 424574
rect 590142 388658 590378 388894
rect 590462 388658 590698 388894
rect 590142 388338 590378 388574
rect 590462 388338 590698 388574
rect 590142 352658 590378 352894
rect 590462 352658 590698 352894
rect 590142 352338 590378 352574
rect 590462 352338 590698 352574
rect 590142 316658 590378 316894
rect 590462 316658 590698 316894
rect 590142 316338 590378 316574
rect 590462 316338 590698 316574
rect 590142 280658 590378 280894
rect 590462 280658 590698 280894
rect 590142 280338 590378 280574
rect 590462 280338 590698 280574
rect 590142 244658 590378 244894
rect 590462 244658 590698 244894
rect 590142 244338 590378 244574
rect 590462 244338 590698 244574
rect 590142 208658 590378 208894
rect 590462 208658 590698 208894
rect 590142 208338 590378 208574
rect 590462 208338 590698 208574
rect 590142 172658 590378 172894
rect 590462 172658 590698 172894
rect 590142 172338 590378 172574
rect 590462 172338 590698 172574
rect 590142 136658 590378 136894
rect 590462 136658 590698 136894
rect 590142 136338 590378 136574
rect 590462 136338 590698 136574
rect 590142 100658 590378 100894
rect 590462 100658 590698 100894
rect 590142 100338 590378 100574
rect 590462 100338 590698 100574
rect 590142 64658 590378 64894
rect 590462 64658 590698 64894
rect 590142 64338 590378 64574
rect 590462 64338 590698 64574
rect 590142 28658 590378 28894
rect 590462 28658 590698 28894
rect 590142 28338 590378 28574
rect 590462 28338 590698 28574
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 698378 591338 698614
rect 591422 698378 591658 698614
rect 591102 698058 591338 698294
rect 591422 698058 591658 698294
rect 591102 662378 591338 662614
rect 591422 662378 591658 662614
rect 591102 662058 591338 662294
rect 591422 662058 591658 662294
rect 591102 626378 591338 626614
rect 591422 626378 591658 626614
rect 591102 626058 591338 626294
rect 591422 626058 591658 626294
rect 591102 590378 591338 590614
rect 591422 590378 591658 590614
rect 591102 590058 591338 590294
rect 591422 590058 591658 590294
rect 591102 554378 591338 554614
rect 591422 554378 591658 554614
rect 591102 554058 591338 554294
rect 591422 554058 591658 554294
rect 591102 518378 591338 518614
rect 591422 518378 591658 518614
rect 591102 518058 591338 518294
rect 591422 518058 591658 518294
rect 591102 482378 591338 482614
rect 591422 482378 591658 482614
rect 591102 482058 591338 482294
rect 591422 482058 591658 482294
rect 591102 446378 591338 446614
rect 591422 446378 591658 446614
rect 591102 446058 591338 446294
rect 591422 446058 591658 446294
rect 591102 410378 591338 410614
rect 591422 410378 591658 410614
rect 591102 410058 591338 410294
rect 591422 410058 591658 410294
rect 591102 374378 591338 374614
rect 591422 374378 591658 374614
rect 591102 374058 591338 374294
rect 591422 374058 591658 374294
rect 591102 338378 591338 338614
rect 591422 338378 591658 338614
rect 591102 338058 591338 338294
rect 591422 338058 591658 338294
rect 591102 302378 591338 302614
rect 591422 302378 591658 302614
rect 591102 302058 591338 302294
rect 591422 302058 591658 302294
rect 591102 266378 591338 266614
rect 591422 266378 591658 266614
rect 591102 266058 591338 266294
rect 591422 266058 591658 266294
rect 591102 230378 591338 230614
rect 591422 230378 591658 230614
rect 591102 230058 591338 230294
rect 591422 230058 591658 230294
rect 591102 194378 591338 194614
rect 591422 194378 591658 194614
rect 591102 194058 591338 194294
rect 591422 194058 591658 194294
rect 591102 158378 591338 158614
rect 591422 158378 591658 158614
rect 591102 158058 591338 158294
rect 591422 158058 591658 158294
rect 591102 122378 591338 122614
rect 591422 122378 591658 122614
rect 591102 122058 591338 122294
rect 591422 122058 591658 122294
rect 591102 86378 591338 86614
rect 591422 86378 591658 86614
rect 591102 86058 591338 86294
rect 591422 86058 591658 86294
rect 591102 50378 591338 50614
rect 591422 50378 591658 50614
rect 591102 50058 591338 50294
rect 591422 50058 591658 50294
rect 591102 14378 591338 14614
rect 591422 14378 591658 14614
rect 591102 14058 591338 14294
rect 591422 14058 591658 14294
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 680378 592298 680614
rect 592382 680378 592618 680614
rect 592062 680058 592298 680294
rect 592382 680058 592618 680294
rect 592062 644378 592298 644614
rect 592382 644378 592618 644614
rect 592062 644058 592298 644294
rect 592382 644058 592618 644294
rect 592062 608378 592298 608614
rect 592382 608378 592618 608614
rect 592062 608058 592298 608294
rect 592382 608058 592618 608294
rect 592062 572378 592298 572614
rect 592382 572378 592618 572614
rect 592062 572058 592298 572294
rect 592382 572058 592618 572294
rect 592062 536378 592298 536614
rect 592382 536378 592618 536614
rect 592062 536058 592298 536294
rect 592382 536058 592618 536294
rect 592062 500378 592298 500614
rect 592382 500378 592618 500614
rect 592062 500058 592298 500294
rect 592382 500058 592618 500294
rect 592062 464378 592298 464614
rect 592382 464378 592618 464614
rect 592062 464058 592298 464294
rect 592382 464058 592618 464294
rect 592062 428378 592298 428614
rect 592382 428378 592618 428614
rect 592062 428058 592298 428294
rect 592382 428058 592618 428294
rect 592062 392378 592298 392614
rect 592382 392378 592618 392614
rect 592062 392058 592298 392294
rect 592382 392058 592618 392294
rect 592062 356378 592298 356614
rect 592382 356378 592618 356614
rect 592062 356058 592298 356294
rect 592382 356058 592618 356294
rect 592062 320378 592298 320614
rect 592382 320378 592618 320614
rect 592062 320058 592298 320294
rect 592382 320058 592618 320294
rect 592062 284378 592298 284614
rect 592382 284378 592618 284614
rect 592062 284058 592298 284294
rect 592382 284058 592618 284294
rect 592062 248378 592298 248614
rect 592382 248378 592618 248614
rect 592062 248058 592298 248294
rect 592382 248058 592618 248294
rect 592062 212378 592298 212614
rect 592382 212378 592618 212614
rect 592062 212058 592298 212294
rect 592382 212058 592618 212294
rect 592062 176378 592298 176614
rect 592382 176378 592618 176614
rect 592062 176058 592298 176294
rect 592382 176058 592618 176294
rect 592062 140378 592298 140614
rect 592382 140378 592618 140614
rect 592062 140058 592298 140294
rect 592382 140058 592618 140294
rect 592062 104378 592298 104614
rect 592382 104378 592618 104614
rect 592062 104058 592298 104294
rect 592382 104058 592618 104294
rect 592062 68378 592298 68614
rect 592382 68378 592618 68614
rect 592062 68058 592298 68294
rect 592382 68058 592618 68294
rect 592062 32378 592298 32614
rect 592382 32378 592618 32614
rect 592062 32058 592298 32294
rect 592382 32058 592618 32294
rect 570986 -7302 571222 -7066
rect 571306 -7302 571542 -7066
rect 570986 -7622 571222 -7386
rect 571306 -7622 571542 -7386
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 592650 698294
rect -8726 698026 592650 698058
rect -6806 694894 590730 694926
rect -6806 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 590730 694894
rect -6806 694574 590730 694658
rect -6806 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 590730 694574
rect -6806 694306 590730 694338
rect -4886 691174 588810 691206
rect -4886 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 588810 691174
rect -4886 690854 588810 690938
rect -4886 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 588810 690854
rect -4886 690586 588810 690618
rect -2966 687454 586890 687486
rect -2966 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 586890 687454
rect -2966 687134 586890 687218
rect -2966 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 586890 687134
rect -2966 686866 586890 686898
rect -8726 680614 592650 680646
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect -8726 680294 592650 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect -8726 680026 592650 680058
rect -6806 676894 590730 676926
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect -6806 676574 590730 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect -6806 676306 590730 676338
rect -4886 673174 588810 673206
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect -4886 672854 588810 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect -4886 672586 588810 672618
rect -2966 669454 586890 669486
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect -2966 669134 586890 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect -2966 668866 586890 668898
rect -8726 662614 592650 662646
rect -8726 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 592650 662294
rect -8726 662026 592650 662058
rect -6806 658894 590730 658926
rect -6806 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 590730 658894
rect -6806 658574 590730 658658
rect -6806 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 590730 658574
rect -6806 658306 590730 658338
rect -4886 655174 588810 655206
rect -4886 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 588810 655174
rect -4886 654854 588810 654938
rect -4886 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 588810 654854
rect -4886 654586 588810 654618
rect -2966 651454 586890 651486
rect -2966 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 586890 651454
rect -2966 651134 586890 651218
rect -2966 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 586890 651134
rect -2966 650866 586890 650898
rect -8726 644614 592650 644646
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect -8726 644294 592650 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect -8726 644026 592650 644058
rect -6806 640894 590730 640926
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect -6806 640574 590730 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect -6806 640306 590730 640338
rect -4886 637174 588810 637206
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect -4886 636854 588810 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect -4886 636586 588810 636618
rect -2966 633454 586890 633486
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect -2966 633134 586890 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect -2966 632866 586890 632898
rect -8726 626614 592650 626646
rect -8726 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 592650 626294
rect -8726 626026 592650 626058
rect -6806 622894 590730 622926
rect -6806 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 590730 622894
rect -6806 622574 590730 622658
rect -6806 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 590730 622574
rect -6806 622306 590730 622338
rect -4886 619174 588810 619206
rect -4886 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 588810 619174
rect -4886 618854 588810 618938
rect -4886 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 588810 618854
rect -4886 618586 588810 618618
rect -2966 615454 586890 615486
rect -2966 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 586890 615454
rect -2966 615134 586890 615218
rect -2966 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 586890 615134
rect -2966 614866 586890 614898
rect -8726 608614 592650 608646
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect -8726 608294 592650 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect -8726 608026 592650 608058
rect -6806 604894 590730 604926
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect -6806 604574 590730 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect -6806 604306 590730 604338
rect -4886 601174 588810 601206
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect -4886 600854 588810 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect -4886 600586 588810 600618
rect -2966 597454 586890 597486
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect -2966 597134 586890 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect -2966 596866 586890 596898
rect -8726 590614 592650 590646
rect -8726 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 592650 590294
rect -8726 590026 592650 590058
rect -6806 586894 590730 586926
rect -6806 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 590730 586894
rect -6806 586574 590730 586658
rect -6806 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 590730 586574
rect -6806 586306 590730 586338
rect -4886 583174 588810 583206
rect -4886 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 77546 583174
rect 77782 582938 77866 583174
rect 78102 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 588810 583174
rect -4886 582854 588810 582938
rect -4886 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 77546 582854
rect 77782 582618 77866 582854
rect 78102 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 588810 582854
rect -4886 582586 588810 582618
rect -2966 579454 586890 579486
rect -2966 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 586890 579454
rect -2966 579134 586890 579218
rect -2966 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 586890 579134
rect -2966 578866 586890 578898
rect -8726 572614 592650 572646
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect -8726 572294 592650 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect -8726 572026 592650 572058
rect -6806 568894 590730 568926
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect -6806 568574 590730 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect -6806 568306 590730 568338
rect -4886 565174 588810 565206
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect -4886 564854 588810 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect -4886 564586 588810 564618
rect -2966 561454 586890 561486
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect -2966 561134 586890 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect -2966 560866 586890 560898
rect -8726 554614 592650 554646
rect -8726 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 84986 554614
rect 85222 554378 85306 554614
rect 85542 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 84986 554294
rect 85222 554058 85306 554294
rect 85542 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 592650 554294
rect -8726 554026 592650 554058
rect -6806 550894 590730 550926
rect -6806 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 81266 550894
rect 81502 550658 81586 550894
rect 81822 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 590730 550894
rect -6806 550574 590730 550658
rect -6806 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 81266 550574
rect 81502 550338 81586 550574
rect 81822 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 590730 550574
rect -6806 550306 590730 550338
rect -4886 547174 588810 547206
rect -4886 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 77546 547174
rect 77782 546938 77866 547174
rect 78102 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 588810 547174
rect -4886 546854 588810 546938
rect -4886 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 77546 546854
rect 77782 546618 77866 546854
rect 78102 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 588810 546854
rect -4886 546586 588810 546618
rect -2966 543454 586890 543486
rect -2966 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 586890 543454
rect -2966 543134 586890 543218
rect -2966 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 586890 543134
rect -2966 542866 586890 542898
rect -8726 536614 592650 536646
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 210986 536614
rect 211222 536378 211306 536614
rect 211542 536378 246986 536614
rect 247222 536378 247306 536614
rect 247542 536378 282986 536614
rect 283222 536378 283306 536614
rect 283542 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 354986 536614
rect 355222 536378 355306 536614
rect 355542 536378 390986 536614
rect 391222 536378 391306 536614
rect 391542 536378 426986 536614
rect 427222 536378 427306 536614
rect 427542 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect -8726 536294 592650 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 210986 536294
rect 211222 536058 211306 536294
rect 211542 536058 246986 536294
rect 247222 536058 247306 536294
rect 247542 536058 282986 536294
rect 283222 536058 283306 536294
rect 283542 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 354986 536294
rect 355222 536058 355306 536294
rect 355542 536058 390986 536294
rect 391222 536058 391306 536294
rect 391542 536058 426986 536294
rect 427222 536058 427306 536294
rect 427542 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect -8726 536026 592650 536058
rect -6806 532894 590730 532926
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 207266 532894
rect 207502 532658 207586 532894
rect 207822 532658 243266 532894
rect 243502 532658 243586 532894
rect 243822 532658 279266 532894
rect 279502 532658 279586 532894
rect 279822 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 351266 532894
rect 351502 532658 351586 532894
rect 351822 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 423266 532894
rect 423502 532658 423586 532894
rect 423822 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect -6806 532574 590730 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 207266 532574
rect 207502 532338 207586 532574
rect 207822 532338 243266 532574
rect 243502 532338 243586 532574
rect 243822 532338 279266 532574
rect 279502 532338 279586 532574
rect 279822 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 351266 532574
rect 351502 532338 351586 532574
rect 351822 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 423266 532574
rect 423502 532338 423586 532574
rect 423822 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect -6806 532306 590730 532338
rect -4886 529174 588810 529206
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 203546 529174
rect 203782 528938 203866 529174
rect 204102 528938 239546 529174
rect 239782 528938 239866 529174
rect 240102 528938 275546 529174
rect 275782 528938 275866 529174
rect 276102 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 347546 529174
rect 347782 528938 347866 529174
rect 348102 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect -4886 528854 588810 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 203546 528854
rect 203782 528618 203866 528854
rect 204102 528618 239546 528854
rect 239782 528618 239866 528854
rect 240102 528618 275546 528854
rect 275782 528618 275866 528854
rect 276102 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 347546 528854
rect 347782 528618 347866 528854
rect 348102 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect -4886 528586 588810 528618
rect -2966 525454 586890 525486
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect -2966 525134 586890 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect -2966 524866 586890 524898
rect -8726 518614 592650 518646
rect -8726 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 592650 518294
rect -8726 518026 592650 518058
rect -6806 514894 590730 514926
rect -6806 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 590730 514894
rect -6806 514574 590730 514658
rect -6806 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 590730 514574
rect -6806 514306 590730 514338
rect -4886 511174 588810 511206
rect -4886 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 588810 511174
rect -4886 510854 588810 510938
rect -4886 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 588810 510854
rect -4886 510586 588810 510618
rect -2966 507454 586890 507486
rect -2966 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 586890 507454
rect -2966 507134 586890 507218
rect -2966 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 586890 507134
rect -2966 506866 586890 506898
rect -8726 500614 592650 500646
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 174986 500614
rect 175222 500378 175306 500614
rect 175542 500378 210986 500614
rect 211222 500378 211306 500614
rect 211542 500378 246986 500614
rect 247222 500378 247306 500614
rect 247542 500378 282986 500614
rect 283222 500378 283306 500614
rect 283542 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect -8726 500294 592650 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 174986 500294
rect 175222 500058 175306 500294
rect 175542 500058 210986 500294
rect 211222 500058 211306 500294
rect 211542 500058 246986 500294
rect 247222 500058 247306 500294
rect 247542 500058 282986 500294
rect 283222 500058 283306 500294
rect 283542 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect -8726 500026 592650 500058
rect -6806 496894 590730 496926
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 171266 496894
rect 171502 496658 171586 496894
rect 171822 496658 207266 496894
rect 207502 496658 207586 496894
rect 207822 496658 243266 496894
rect 243502 496658 243586 496894
rect 243822 496658 279266 496894
rect 279502 496658 279586 496894
rect 279822 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect -6806 496574 590730 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 171266 496574
rect 171502 496338 171586 496574
rect 171822 496338 207266 496574
rect 207502 496338 207586 496574
rect 207822 496338 243266 496574
rect 243502 496338 243586 496574
rect 243822 496338 279266 496574
rect 279502 496338 279586 496574
rect 279822 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect -6806 496306 590730 496338
rect -4886 493174 588810 493206
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 167546 493174
rect 167782 492938 167866 493174
rect 168102 492938 203546 493174
rect 203782 492938 203866 493174
rect 204102 492938 239546 493174
rect 239782 492938 239866 493174
rect 240102 492938 275546 493174
rect 275782 492938 275866 493174
rect 276102 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect -4886 492854 588810 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 167546 492854
rect 167782 492618 167866 492854
rect 168102 492618 203546 492854
rect 203782 492618 203866 492854
rect 204102 492618 239546 492854
rect 239782 492618 239866 492854
rect 240102 492618 275546 492854
rect 275782 492618 275866 492854
rect 276102 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect -4886 492586 588810 492618
rect -2966 489454 586890 489486
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect -2966 489134 586890 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect -2966 488866 586890 488898
rect -8726 482614 592650 482646
rect -8726 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 592650 482294
rect -8726 482026 592650 482058
rect -6806 478894 590730 478926
rect -6806 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 590730 478894
rect -6806 478574 590730 478658
rect -6806 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 590730 478574
rect -6806 478306 590730 478338
rect -4886 475174 588810 475206
rect -4886 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 588810 475174
rect -4886 474854 588810 474938
rect -4886 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 588810 474854
rect -4886 474586 588810 474618
rect -2966 471454 586890 471486
rect -2966 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 586890 471454
rect -2966 471134 586890 471218
rect -2966 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 586890 471134
rect -2966 470866 586890 470898
rect -8726 464614 592650 464646
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 246986 464614
rect 247222 464378 247306 464614
rect 247542 464378 282986 464614
rect 283222 464378 283306 464614
rect 283542 464378 318986 464614
rect 319222 464378 319306 464614
rect 319542 464378 354986 464614
rect 355222 464378 355306 464614
rect 355542 464378 390986 464614
rect 391222 464378 391306 464614
rect 391542 464378 426986 464614
rect 427222 464378 427306 464614
rect 427542 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect -8726 464294 592650 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 246986 464294
rect 247222 464058 247306 464294
rect 247542 464058 282986 464294
rect 283222 464058 283306 464294
rect 283542 464058 318986 464294
rect 319222 464058 319306 464294
rect 319542 464058 354986 464294
rect 355222 464058 355306 464294
rect 355542 464058 390986 464294
rect 391222 464058 391306 464294
rect 391542 464058 426986 464294
rect 427222 464058 427306 464294
rect 427542 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect -8726 464026 592650 464058
rect -6806 460894 590730 460926
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 243266 460894
rect 243502 460658 243586 460894
rect 243822 460658 279266 460894
rect 279502 460658 279586 460894
rect 279822 460658 315266 460894
rect 315502 460658 315586 460894
rect 315822 460658 351266 460894
rect 351502 460658 351586 460894
rect 351822 460658 387266 460894
rect 387502 460658 387586 460894
rect 387822 460658 423266 460894
rect 423502 460658 423586 460894
rect 423822 460658 459266 460894
rect 459502 460658 459586 460894
rect 459822 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect -6806 460574 590730 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 243266 460574
rect 243502 460338 243586 460574
rect 243822 460338 279266 460574
rect 279502 460338 279586 460574
rect 279822 460338 315266 460574
rect 315502 460338 315586 460574
rect 315822 460338 351266 460574
rect 351502 460338 351586 460574
rect 351822 460338 387266 460574
rect 387502 460338 387586 460574
rect 387822 460338 423266 460574
rect 423502 460338 423586 460574
rect 423822 460338 459266 460574
rect 459502 460338 459586 460574
rect 459822 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect -6806 460306 590730 460338
rect -4886 457174 588810 457206
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 239546 457174
rect 239782 456938 239866 457174
rect 240102 456938 275546 457174
rect 275782 456938 275866 457174
rect 276102 456938 311546 457174
rect 311782 456938 311866 457174
rect 312102 456938 347546 457174
rect 347782 456938 347866 457174
rect 348102 456938 383546 457174
rect 383782 456938 383866 457174
rect 384102 456938 419546 457174
rect 419782 456938 419866 457174
rect 420102 456938 455546 457174
rect 455782 456938 455866 457174
rect 456102 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect -4886 456854 588810 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 239546 456854
rect 239782 456618 239866 456854
rect 240102 456618 275546 456854
rect 275782 456618 275866 456854
rect 276102 456618 311546 456854
rect 311782 456618 311866 456854
rect 312102 456618 347546 456854
rect 347782 456618 347866 456854
rect 348102 456618 383546 456854
rect 383782 456618 383866 456854
rect 384102 456618 419546 456854
rect 419782 456618 419866 456854
rect 420102 456618 455546 456854
rect 455782 456618 455866 456854
rect 456102 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect -4886 456586 588810 456618
rect -2966 453454 586890 453486
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 50328 453454
rect 50564 453218 186056 453454
rect 186292 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect -2966 453134 586890 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 50328 453134
rect 50564 452898 186056 453134
rect 186292 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect -2966 452866 586890 452898
rect -8726 446614 592650 446646
rect -8726 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 192986 446614
rect 193222 446378 193306 446614
rect 193542 446378 228986 446614
rect 229222 446378 229306 446614
rect 229542 446378 264986 446614
rect 265222 446378 265306 446614
rect 265542 446378 300986 446614
rect 301222 446378 301306 446614
rect 301542 446378 336986 446614
rect 337222 446378 337306 446614
rect 337542 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 192986 446294
rect 193222 446058 193306 446294
rect 193542 446058 228986 446294
rect 229222 446058 229306 446294
rect 229542 446058 264986 446294
rect 265222 446058 265306 446294
rect 265542 446058 300986 446294
rect 301222 446058 301306 446294
rect 301542 446058 336986 446294
rect 337222 446058 337306 446294
rect 337542 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 592650 446294
rect -8726 446026 592650 446058
rect -6806 442894 590730 442926
rect -6806 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 225266 442894
rect 225502 442658 225586 442894
rect 225822 442658 261266 442894
rect 261502 442658 261586 442894
rect 261822 442658 297266 442894
rect 297502 442658 297586 442894
rect 297822 442658 333266 442894
rect 333502 442658 333586 442894
rect 333822 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 441266 442894
rect 441502 442658 441586 442894
rect 441822 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 590730 442894
rect -6806 442574 590730 442658
rect -6806 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 225266 442574
rect 225502 442338 225586 442574
rect 225822 442338 261266 442574
rect 261502 442338 261586 442574
rect 261822 442338 297266 442574
rect 297502 442338 297586 442574
rect 297822 442338 333266 442574
rect 333502 442338 333586 442574
rect 333822 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 441266 442574
rect 441502 442338 441586 442574
rect 441822 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 590730 442574
rect -6806 442306 590730 442338
rect -4886 439174 588810 439206
rect -4886 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 221546 439174
rect 221782 438938 221866 439174
rect 222102 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 588810 439174
rect -4886 438854 588810 438938
rect -4886 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 221546 438854
rect 221782 438618 221866 438854
rect 222102 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 588810 438854
rect -4886 438586 588810 438618
rect -2966 435454 586890 435486
rect -2966 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 51008 435454
rect 51244 435218 185376 435454
rect 185612 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 244250 435454
rect 244486 435218 274970 435454
rect 275206 435218 305690 435454
rect 305926 435218 336410 435454
rect 336646 435218 367130 435454
rect 367366 435218 397850 435454
rect 398086 435218 428570 435454
rect 428806 435218 459290 435454
rect 459526 435218 490010 435454
rect 490246 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 586890 435454
rect -2966 435134 586890 435218
rect -2966 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 51008 435134
rect 51244 434898 185376 435134
rect 185612 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 244250 435134
rect 244486 434898 274970 435134
rect 275206 434898 305690 435134
rect 305926 434898 336410 435134
rect 336646 434898 367130 435134
rect 367366 434898 397850 435134
rect 398086 434898 428570 435134
rect 428806 434898 459290 435134
rect 459526 434898 490010 435134
rect 490246 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 586890 435134
rect -2966 434866 586890 434898
rect -8726 428614 592650 428646
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 210986 428614
rect 211222 428378 211306 428614
rect 211542 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect -8726 428294 592650 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 210986 428294
rect 211222 428058 211306 428294
rect 211542 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect -8726 428026 592650 428058
rect -6806 424894 590730 424926
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 207266 424894
rect 207502 424658 207586 424894
rect 207822 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect -6806 424574 590730 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 207266 424574
rect 207502 424338 207586 424574
rect 207822 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect -6806 424306 590730 424338
rect -4886 421174 588810 421206
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 203546 421174
rect 203782 420938 203866 421174
rect 204102 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect -4886 420854 588810 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 203546 420854
rect 203782 420618 203866 420854
rect 204102 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect -4886 420586 588810 420618
rect -2966 417454 586890 417486
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 50328 417454
rect 50564 417218 186056 417454
rect 186292 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 259610 417454
rect 259846 417218 290330 417454
rect 290566 417218 321050 417454
rect 321286 417218 351770 417454
rect 352006 417218 382490 417454
rect 382726 417218 413210 417454
rect 413446 417218 443930 417454
rect 444166 417218 474650 417454
rect 474886 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect -2966 417134 586890 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 50328 417134
rect 50564 416898 186056 417134
rect 186292 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 259610 417134
rect 259846 416898 290330 417134
rect 290566 416898 321050 417134
rect 321286 416898 351770 417134
rect 352006 416898 382490 417134
rect 382726 416898 413210 417134
rect 413446 416898 443930 417134
rect 444166 416898 474650 417134
rect 474886 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect -2966 416866 586890 416898
rect -8726 410614 592650 410646
rect -8726 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 192986 410614
rect 193222 410378 193306 410614
rect 193542 410378 228986 410614
rect 229222 410378 229306 410614
rect 229542 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 192986 410294
rect 193222 410058 193306 410294
rect 193542 410058 228986 410294
rect 229222 410058 229306 410294
rect 229542 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 592650 410294
rect -8726 410026 592650 410058
rect -6806 406894 590730 406926
rect -6806 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 189266 406894
rect 189502 406658 189586 406894
rect 189822 406658 225266 406894
rect 225502 406658 225586 406894
rect 225822 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 590730 406894
rect -6806 406574 590730 406658
rect -6806 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 189266 406574
rect 189502 406338 189586 406574
rect 189822 406338 225266 406574
rect 225502 406338 225586 406574
rect 225822 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 590730 406574
rect -6806 406306 590730 406338
rect -4886 403174 588810 403206
rect -4886 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 221546 403174
rect 221782 402938 221866 403174
rect 222102 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 588810 403174
rect -4886 402854 588810 402938
rect -4886 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 221546 402854
rect 221782 402618 221866 402854
rect 222102 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 588810 402854
rect -4886 402586 588810 402618
rect -2966 399454 586890 399486
rect -2966 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 51008 399454
rect 51244 399218 185376 399454
rect 185612 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 244250 399454
rect 244486 399218 274970 399454
rect 275206 399218 305690 399454
rect 305926 399218 336410 399454
rect 336646 399218 367130 399454
rect 367366 399218 397850 399454
rect 398086 399218 428570 399454
rect 428806 399218 459290 399454
rect 459526 399218 490010 399454
rect 490246 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 586890 399454
rect -2966 399134 586890 399218
rect -2966 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 51008 399134
rect 51244 398898 185376 399134
rect 185612 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 244250 399134
rect 244486 398898 274970 399134
rect 275206 398898 305690 399134
rect 305926 398898 336410 399134
rect 336646 398898 367130 399134
rect 367366 398898 397850 399134
rect 398086 398898 428570 399134
rect 428806 398898 459290 399134
rect 459526 398898 490010 399134
rect 490246 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 586890 399134
rect -2966 398866 586890 398898
rect -8726 392614 592650 392646
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 210986 392614
rect 211222 392378 211306 392614
rect 211542 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect -8726 392294 592650 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 210986 392294
rect 211222 392058 211306 392294
rect 211542 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect -8726 392026 592650 392058
rect -6806 388894 590730 388926
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 207266 388894
rect 207502 388658 207586 388894
rect 207822 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect -6806 388574 590730 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 207266 388574
rect 207502 388338 207586 388574
rect 207822 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect -6806 388306 590730 388338
rect -4886 385174 588810 385206
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 203546 385174
rect 203782 384938 203866 385174
rect 204102 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect -4886 384854 588810 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 203546 384854
rect 203782 384618 203866 384854
rect 204102 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect -4886 384586 588810 384618
rect -2966 381454 586890 381486
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 50328 381454
rect 50564 381218 186056 381454
rect 186292 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 259610 381454
rect 259846 381218 290330 381454
rect 290566 381218 321050 381454
rect 321286 381218 351770 381454
rect 352006 381218 382490 381454
rect 382726 381218 413210 381454
rect 413446 381218 443930 381454
rect 444166 381218 474650 381454
rect 474886 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect -2966 381134 586890 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 50328 381134
rect 50564 380898 186056 381134
rect 186292 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 259610 381134
rect 259846 380898 290330 381134
rect 290566 380898 321050 381134
rect 321286 380898 351770 381134
rect 352006 380898 382490 381134
rect 382726 380898 413210 381134
rect 413446 380898 443930 381134
rect 444166 380898 474650 381134
rect 474886 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect -2966 380866 586890 380898
rect -8726 374614 592650 374646
rect -8726 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 592650 374294
rect -8726 374026 592650 374058
rect -6806 370894 590730 370926
rect -6806 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 590730 370894
rect -6806 370574 590730 370658
rect -6806 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 590730 370574
rect -6806 370306 590730 370338
rect -4886 367174 588810 367206
rect -4886 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 588810 367174
rect -4886 366854 588810 366938
rect -4886 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 588810 366854
rect -4886 366586 588810 366618
rect -2966 363454 586890 363486
rect -2966 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 244250 363454
rect 244486 363218 274970 363454
rect 275206 363218 305690 363454
rect 305926 363218 336410 363454
rect 336646 363218 367130 363454
rect 367366 363218 397850 363454
rect 398086 363218 428570 363454
rect 428806 363218 459290 363454
rect 459526 363218 490010 363454
rect 490246 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 586890 363454
rect -2966 363134 586890 363218
rect -2966 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 244250 363134
rect 244486 362898 274970 363134
rect 275206 362898 305690 363134
rect 305926 362898 336410 363134
rect 336646 362898 367130 363134
rect 367366 362898 397850 363134
rect 398086 362898 428570 363134
rect 428806 362898 459290 363134
rect 459526 362898 490010 363134
rect 490246 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 586890 363134
rect -2966 362866 586890 362898
rect -8726 356614 592650 356646
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 102986 356614
rect 103222 356378 103306 356614
rect 103542 356378 138986 356614
rect 139222 356378 139306 356614
rect 139542 356378 174986 356614
rect 175222 356378 175306 356614
rect 175542 356378 210986 356614
rect 211222 356378 211306 356614
rect 211542 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect -8726 356294 592650 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 102986 356294
rect 103222 356058 103306 356294
rect 103542 356058 138986 356294
rect 139222 356058 139306 356294
rect 139542 356058 174986 356294
rect 175222 356058 175306 356294
rect 175542 356058 210986 356294
rect 211222 356058 211306 356294
rect 211542 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect -8726 356026 592650 356058
rect -6806 352894 590730 352926
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 63266 352894
rect 63502 352658 63586 352894
rect 63822 352658 99266 352894
rect 99502 352658 99586 352894
rect 99822 352658 135266 352894
rect 135502 352658 135586 352894
rect 135822 352658 171266 352894
rect 171502 352658 171586 352894
rect 171822 352658 207266 352894
rect 207502 352658 207586 352894
rect 207822 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect -6806 352574 590730 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 63266 352574
rect 63502 352338 63586 352574
rect 63822 352338 99266 352574
rect 99502 352338 99586 352574
rect 99822 352338 135266 352574
rect 135502 352338 135586 352574
rect 135822 352338 171266 352574
rect 171502 352338 171586 352574
rect 171822 352338 207266 352574
rect 207502 352338 207586 352574
rect 207822 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect -6806 352306 590730 352338
rect -4886 349174 588810 349206
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 59546 349174
rect 59782 348938 59866 349174
rect 60102 348938 95546 349174
rect 95782 348938 95866 349174
rect 96102 348938 131546 349174
rect 131782 348938 131866 349174
rect 132102 348938 167546 349174
rect 167782 348938 167866 349174
rect 168102 348938 203546 349174
rect 203782 348938 203866 349174
rect 204102 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect -4886 348854 588810 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 59546 348854
rect 59782 348618 59866 348854
rect 60102 348618 95546 348854
rect 95782 348618 95866 348854
rect 96102 348618 131546 348854
rect 131782 348618 131866 348854
rect 132102 348618 167546 348854
rect 167782 348618 167866 348854
rect 168102 348618 203546 348854
rect 203782 348618 203866 348854
rect 204102 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect -4886 348586 588810 348618
rect -2966 345454 586890 345486
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 259610 345454
rect 259846 345218 290330 345454
rect 290566 345218 321050 345454
rect 321286 345218 351770 345454
rect 352006 345218 382490 345454
rect 382726 345218 413210 345454
rect 413446 345218 443930 345454
rect 444166 345218 474650 345454
rect 474886 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect -2966 345134 586890 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 259610 345134
rect 259846 344898 290330 345134
rect 290566 344898 321050 345134
rect 321286 344898 351770 345134
rect 352006 344898 382490 345134
rect 382726 344898 413210 345134
rect 413446 344898 443930 345134
rect 444166 344898 474650 345134
rect 474886 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect -2966 344866 586890 344898
rect -8726 338614 592650 338646
rect -8726 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 84986 338614
rect 85222 338378 85306 338614
rect 85542 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 192986 338614
rect 193222 338378 193306 338614
rect 193542 338378 228986 338614
rect 229222 338378 229306 338614
rect 229542 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 84986 338294
rect 85222 338058 85306 338294
rect 85542 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 192986 338294
rect 193222 338058 193306 338294
rect 193542 338058 228986 338294
rect 229222 338058 229306 338294
rect 229542 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 592650 338294
rect -8726 338026 592650 338058
rect -6806 334894 590730 334926
rect -6806 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 189266 334894
rect 189502 334658 189586 334894
rect 189822 334658 225266 334894
rect 225502 334658 225586 334894
rect 225822 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 590730 334894
rect -6806 334574 590730 334658
rect -6806 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 189266 334574
rect 189502 334338 189586 334574
rect 189822 334338 225266 334574
rect 225502 334338 225586 334574
rect 225822 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 590730 334574
rect -6806 334306 590730 334338
rect -4886 331174 588810 331206
rect -4886 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 113546 331174
rect 113782 330938 113866 331174
rect 114102 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 221546 331174
rect 221782 330938 221866 331174
rect 222102 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 588810 331174
rect -4886 330854 588810 330938
rect -4886 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 113546 330854
rect 113782 330618 113866 330854
rect 114102 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 221546 330854
rect 221782 330618 221866 330854
rect 222102 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 588810 330854
rect -4886 330586 588810 330618
rect -2966 327454 586890 327486
rect -2966 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 244250 327454
rect 244486 327218 274970 327454
rect 275206 327218 305690 327454
rect 305926 327218 336410 327454
rect 336646 327218 367130 327454
rect 367366 327218 397850 327454
rect 398086 327218 428570 327454
rect 428806 327218 459290 327454
rect 459526 327218 490010 327454
rect 490246 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 586890 327454
rect -2966 327134 586890 327218
rect -2966 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 244250 327134
rect 244486 326898 274970 327134
rect 275206 326898 305690 327134
rect 305926 326898 336410 327134
rect 336646 326898 367130 327134
rect 367366 326898 397850 327134
rect 398086 326898 428570 327134
rect 428806 326898 459290 327134
rect 459526 326898 490010 327134
rect 490246 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 586890 327134
rect -2966 326866 586890 326898
rect -8726 320614 592650 320646
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 66986 320614
rect 67222 320378 67306 320614
rect 67542 320378 102986 320614
rect 103222 320378 103306 320614
rect 103542 320378 138986 320614
rect 139222 320378 139306 320614
rect 139542 320378 174986 320614
rect 175222 320378 175306 320614
rect 175542 320378 210986 320614
rect 211222 320378 211306 320614
rect 211542 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect -8726 320294 592650 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 66986 320294
rect 67222 320058 67306 320294
rect 67542 320058 102986 320294
rect 103222 320058 103306 320294
rect 103542 320058 138986 320294
rect 139222 320058 139306 320294
rect 139542 320058 174986 320294
rect 175222 320058 175306 320294
rect 175542 320058 210986 320294
rect 211222 320058 211306 320294
rect 211542 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect -8726 320026 592650 320058
rect -6806 316894 590730 316926
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 63266 316894
rect 63502 316658 63586 316894
rect 63822 316658 99266 316894
rect 99502 316658 99586 316894
rect 99822 316658 135266 316894
rect 135502 316658 135586 316894
rect 135822 316658 171266 316894
rect 171502 316658 171586 316894
rect 171822 316658 207266 316894
rect 207502 316658 207586 316894
rect 207822 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect -6806 316574 590730 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 63266 316574
rect 63502 316338 63586 316574
rect 63822 316338 99266 316574
rect 99502 316338 99586 316574
rect 99822 316338 135266 316574
rect 135502 316338 135586 316574
rect 135822 316338 171266 316574
rect 171502 316338 171586 316574
rect 171822 316338 207266 316574
rect 207502 316338 207586 316574
rect 207822 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect -6806 316306 590730 316338
rect -4886 313174 588810 313206
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 59546 313174
rect 59782 312938 59866 313174
rect 60102 312938 95546 313174
rect 95782 312938 95866 313174
rect 96102 312938 131546 313174
rect 131782 312938 131866 313174
rect 132102 312938 167546 313174
rect 167782 312938 167866 313174
rect 168102 312938 203546 313174
rect 203782 312938 203866 313174
rect 204102 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect -4886 312854 588810 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 59546 312854
rect 59782 312618 59866 312854
rect 60102 312618 95546 312854
rect 95782 312618 95866 312854
rect 96102 312618 131546 312854
rect 131782 312618 131866 312854
rect 132102 312618 167546 312854
rect 167782 312618 167866 312854
rect 168102 312618 203546 312854
rect 203782 312618 203866 312854
rect 204102 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect -4886 312586 588810 312618
rect -2966 309454 586890 309486
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 259610 309454
rect 259846 309218 290330 309454
rect 290566 309218 321050 309454
rect 321286 309218 351770 309454
rect 352006 309218 382490 309454
rect 382726 309218 413210 309454
rect 413446 309218 443930 309454
rect 444166 309218 474650 309454
rect 474886 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect -2966 309134 586890 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 259610 309134
rect 259846 308898 290330 309134
rect 290566 308898 321050 309134
rect 321286 308898 351770 309134
rect 352006 308898 382490 309134
rect 382726 308898 413210 309134
rect 413446 308898 443930 309134
rect 444166 308898 474650 309134
rect 474886 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect -2966 308866 586890 308898
rect -8726 302614 592650 302646
rect -8726 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 84986 302614
rect 85222 302378 85306 302614
rect 85542 302378 120986 302614
rect 121222 302378 121306 302614
rect 121542 302378 156986 302614
rect 157222 302378 157306 302614
rect 157542 302378 192986 302614
rect 193222 302378 193306 302614
rect 193542 302378 228986 302614
rect 229222 302378 229306 302614
rect 229542 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 84986 302294
rect 85222 302058 85306 302294
rect 85542 302058 120986 302294
rect 121222 302058 121306 302294
rect 121542 302058 156986 302294
rect 157222 302058 157306 302294
rect 157542 302058 192986 302294
rect 193222 302058 193306 302294
rect 193542 302058 228986 302294
rect 229222 302058 229306 302294
rect 229542 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 592650 302294
rect -8726 302026 592650 302058
rect -6806 298894 590730 298926
rect -6806 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 81266 298894
rect 81502 298658 81586 298894
rect 81822 298658 117266 298894
rect 117502 298658 117586 298894
rect 117822 298658 153266 298894
rect 153502 298658 153586 298894
rect 153822 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 225266 298894
rect 225502 298658 225586 298894
rect 225822 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 590730 298894
rect -6806 298574 590730 298658
rect -6806 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 81266 298574
rect 81502 298338 81586 298574
rect 81822 298338 117266 298574
rect 117502 298338 117586 298574
rect 117822 298338 153266 298574
rect 153502 298338 153586 298574
rect 153822 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 225266 298574
rect 225502 298338 225586 298574
rect 225822 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 590730 298574
rect -6806 298306 590730 298338
rect -4886 295174 588810 295206
rect -4886 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 77546 295174
rect 77782 294938 77866 295174
rect 78102 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 149546 295174
rect 149782 294938 149866 295174
rect 150102 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 221546 295174
rect 221782 294938 221866 295174
rect 222102 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 588810 295174
rect -4886 294854 588810 294938
rect -4886 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 77546 294854
rect 77782 294618 77866 294854
rect 78102 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 149546 294854
rect 149782 294618 149866 294854
rect 150102 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 221546 294854
rect 221782 294618 221866 294854
rect 222102 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 588810 294854
rect -4886 294586 588810 294618
rect -2966 291454 586890 291486
rect -2966 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 244250 291454
rect 244486 291218 274970 291454
rect 275206 291218 305690 291454
rect 305926 291218 336410 291454
rect 336646 291218 367130 291454
rect 367366 291218 397850 291454
rect 398086 291218 428570 291454
rect 428806 291218 459290 291454
rect 459526 291218 490010 291454
rect 490246 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 586890 291454
rect -2966 291134 586890 291218
rect -2966 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 244250 291134
rect 244486 290898 274970 291134
rect 275206 290898 305690 291134
rect 305926 290898 336410 291134
rect 336646 290898 367130 291134
rect 367366 290898 397850 291134
rect 398086 290898 428570 291134
rect 428806 290898 459290 291134
rect 459526 290898 490010 291134
rect 490246 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 586890 291134
rect -2966 290866 586890 290898
rect -8726 284614 592650 284646
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 210986 284614
rect 211222 284378 211306 284614
rect 211542 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect -8726 284294 592650 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 210986 284294
rect 211222 284058 211306 284294
rect 211542 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect -8726 284026 592650 284058
rect -6806 280894 590730 280926
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 207266 280894
rect 207502 280658 207586 280894
rect 207822 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect -6806 280574 590730 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 207266 280574
rect 207502 280338 207586 280574
rect 207822 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect -6806 280306 590730 280338
rect -4886 277174 588810 277206
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 203546 277174
rect 203782 276938 203866 277174
rect 204102 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect -4886 276854 588810 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 203546 276854
rect 203782 276618 203866 276854
rect 204102 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect -4886 276586 588810 276618
rect -2966 273454 586890 273486
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 50328 273454
rect 50564 273218 186056 273454
rect 186292 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 259610 273454
rect 259846 273218 290330 273454
rect 290566 273218 321050 273454
rect 321286 273218 351770 273454
rect 352006 273218 382490 273454
rect 382726 273218 413210 273454
rect 413446 273218 443930 273454
rect 444166 273218 474650 273454
rect 474886 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect -2966 273134 586890 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 50328 273134
rect 50564 272898 186056 273134
rect 186292 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 259610 273134
rect 259846 272898 290330 273134
rect 290566 272898 321050 273134
rect 321286 272898 351770 273134
rect 352006 272898 382490 273134
rect 382726 272898 413210 273134
rect 413446 272898 443930 273134
rect 444166 272898 474650 273134
rect 474886 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect -2966 272866 586890 272898
rect -8726 266614 592650 266646
rect -8726 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 192986 266614
rect 193222 266378 193306 266614
rect 193542 266378 228986 266614
rect 229222 266378 229306 266614
rect 229542 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 192986 266294
rect 193222 266058 193306 266294
rect 193542 266058 228986 266294
rect 229222 266058 229306 266294
rect 229542 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 592650 266294
rect -8726 266026 592650 266058
rect -6806 262894 590730 262926
rect -6806 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 225266 262894
rect 225502 262658 225586 262894
rect 225822 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 590730 262894
rect -6806 262574 590730 262658
rect -6806 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 225266 262574
rect 225502 262338 225586 262574
rect 225822 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 590730 262574
rect -6806 262306 590730 262338
rect -4886 259174 588810 259206
rect -4886 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 221546 259174
rect 221782 258938 221866 259174
rect 222102 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 588810 259174
rect -4886 258854 588810 258938
rect -4886 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 221546 258854
rect 221782 258618 221866 258854
rect 222102 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 588810 258854
rect -4886 258586 588810 258618
rect -2966 255454 586890 255486
rect -2966 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 51008 255454
rect 51244 255218 185376 255454
rect 185612 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 244250 255454
rect 244486 255218 274970 255454
rect 275206 255218 305690 255454
rect 305926 255218 336410 255454
rect 336646 255218 367130 255454
rect 367366 255218 397850 255454
rect 398086 255218 428570 255454
rect 428806 255218 459290 255454
rect 459526 255218 490010 255454
rect 490246 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 586890 255454
rect -2966 255134 586890 255218
rect -2966 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 51008 255134
rect 51244 254898 185376 255134
rect 185612 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 244250 255134
rect 244486 254898 274970 255134
rect 275206 254898 305690 255134
rect 305926 254898 336410 255134
rect 336646 254898 367130 255134
rect 367366 254898 397850 255134
rect 398086 254898 428570 255134
rect 428806 254898 459290 255134
rect 459526 254898 490010 255134
rect 490246 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 586890 255134
rect -2966 254866 586890 254898
rect -8726 248614 592650 248646
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 210986 248614
rect 211222 248378 211306 248614
rect 211542 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect -8726 248294 592650 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 210986 248294
rect 211222 248058 211306 248294
rect 211542 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect -8726 248026 592650 248058
rect -6806 244894 590730 244926
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 207266 244894
rect 207502 244658 207586 244894
rect 207822 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect -6806 244574 590730 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 207266 244574
rect 207502 244338 207586 244574
rect 207822 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect -6806 244306 590730 244338
rect -4886 241174 588810 241206
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 203546 241174
rect 203782 240938 203866 241174
rect 204102 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect -4886 240854 588810 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 203546 240854
rect 203782 240618 203866 240854
rect 204102 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect -4886 240586 588810 240618
rect -2966 237454 586890 237486
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 50328 237454
rect 50564 237218 186056 237454
rect 186292 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 259610 237454
rect 259846 237218 290330 237454
rect 290566 237218 321050 237454
rect 321286 237218 351770 237454
rect 352006 237218 382490 237454
rect 382726 237218 413210 237454
rect 413446 237218 443930 237454
rect 444166 237218 474650 237454
rect 474886 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect -2966 237134 586890 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 50328 237134
rect 50564 236898 186056 237134
rect 186292 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 259610 237134
rect 259846 236898 290330 237134
rect 290566 236898 321050 237134
rect 321286 236898 351770 237134
rect 352006 236898 382490 237134
rect 382726 236898 413210 237134
rect 413446 236898 443930 237134
rect 444166 236898 474650 237134
rect 474886 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect -2966 236866 586890 236898
rect -8726 230614 592650 230646
rect -8726 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 192986 230614
rect 193222 230378 193306 230614
rect 193542 230378 228986 230614
rect 229222 230378 229306 230614
rect 229542 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 192986 230294
rect 193222 230058 193306 230294
rect 193542 230058 228986 230294
rect 229222 230058 229306 230294
rect 229542 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 592650 230294
rect -8726 230026 592650 230058
rect -6806 226894 590730 226926
rect -6806 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 189266 226894
rect 189502 226658 189586 226894
rect 189822 226658 225266 226894
rect 225502 226658 225586 226894
rect 225822 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 590730 226894
rect -6806 226574 590730 226658
rect -6806 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 189266 226574
rect 189502 226338 189586 226574
rect 189822 226338 225266 226574
rect 225502 226338 225586 226574
rect 225822 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 590730 226574
rect -6806 226306 590730 226338
rect -4886 223174 588810 223206
rect -4886 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 221546 223174
rect 221782 222938 221866 223174
rect 222102 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 588810 223174
rect -4886 222854 588810 222938
rect -4886 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 221546 222854
rect 221782 222618 221866 222854
rect 222102 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 588810 222854
rect -4886 222586 588810 222618
rect -2966 219454 586890 219486
rect -2966 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 51008 219454
rect 51244 219218 185376 219454
rect 185612 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 244250 219454
rect 244486 219218 274970 219454
rect 275206 219218 305690 219454
rect 305926 219218 336410 219454
rect 336646 219218 367130 219454
rect 367366 219218 397850 219454
rect 398086 219218 428570 219454
rect 428806 219218 459290 219454
rect 459526 219218 490010 219454
rect 490246 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 586890 219454
rect -2966 219134 586890 219218
rect -2966 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 51008 219134
rect 51244 218898 185376 219134
rect 185612 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 244250 219134
rect 244486 218898 274970 219134
rect 275206 218898 305690 219134
rect 305926 218898 336410 219134
rect 336646 218898 367130 219134
rect 367366 218898 397850 219134
rect 398086 218898 428570 219134
rect 428806 218898 459290 219134
rect 459526 218898 490010 219134
rect 490246 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 586890 219134
rect -2966 218866 586890 218898
rect -8726 212614 592650 212646
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 210986 212614
rect 211222 212378 211306 212614
rect 211542 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect -8726 212294 592650 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 210986 212294
rect 211222 212058 211306 212294
rect 211542 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect -8726 212026 592650 212058
rect -6806 208894 590730 208926
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 207266 208894
rect 207502 208658 207586 208894
rect 207822 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect -6806 208574 590730 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 207266 208574
rect 207502 208338 207586 208574
rect 207822 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect -6806 208306 590730 208338
rect -4886 205174 588810 205206
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 203546 205174
rect 203782 204938 203866 205174
rect 204102 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect -4886 204854 588810 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 203546 204854
rect 203782 204618 203866 204854
rect 204102 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect -4886 204586 588810 204618
rect -2966 201454 586890 201486
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 50328 201454
rect 50564 201218 186056 201454
rect 186292 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 259610 201454
rect 259846 201218 290330 201454
rect 290566 201218 321050 201454
rect 321286 201218 351770 201454
rect 352006 201218 382490 201454
rect 382726 201218 413210 201454
rect 413446 201218 443930 201454
rect 444166 201218 474650 201454
rect 474886 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect -2966 201134 586890 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 50328 201134
rect 50564 200898 186056 201134
rect 186292 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 259610 201134
rect 259846 200898 290330 201134
rect 290566 200898 321050 201134
rect 321286 200898 351770 201134
rect 352006 200898 382490 201134
rect 382726 200898 413210 201134
rect 413446 200898 443930 201134
rect 444166 200898 474650 201134
rect 474886 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect -2966 200866 586890 200898
rect -8726 194614 592650 194646
rect -8726 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 120986 194614
rect 121222 194378 121306 194614
rect 121542 194378 156986 194614
rect 157222 194378 157306 194614
rect 157542 194378 192986 194614
rect 193222 194378 193306 194614
rect 193542 194378 228986 194614
rect 229222 194378 229306 194614
rect 229542 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 120986 194294
rect 121222 194058 121306 194294
rect 121542 194058 156986 194294
rect 157222 194058 157306 194294
rect 157542 194058 192986 194294
rect 193222 194058 193306 194294
rect 193542 194058 228986 194294
rect 229222 194058 229306 194294
rect 229542 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 592650 194294
rect -8726 194026 592650 194058
rect -6806 190894 590730 190926
rect -6806 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 117266 190894
rect 117502 190658 117586 190894
rect 117822 190658 153266 190894
rect 153502 190658 153586 190894
rect 153822 190658 189266 190894
rect 189502 190658 189586 190894
rect 189822 190658 225266 190894
rect 225502 190658 225586 190894
rect 225822 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 590730 190894
rect -6806 190574 590730 190658
rect -6806 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 117266 190574
rect 117502 190338 117586 190574
rect 117822 190338 153266 190574
rect 153502 190338 153586 190574
rect 153822 190338 189266 190574
rect 189502 190338 189586 190574
rect 189822 190338 225266 190574
rect 225502 190338 225586 190574
rect 225822 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 590730 190574
rect -6806 190306 590730 190338
rect -4886 187174 588810 187206
rect -4886 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 149546 187174
rect 149782 186938 149866 187174
rect 150102 186938 185546 187174
rect 185782 186938 185866 187174
rect 186102 186938 221546 187174
rect 221782 186938 221866 187174
rect 222102 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 588810 187174
rect -4886 186854 588810 186938
rect -4886 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 149546 186854
rect 149782 186618 149866 186854
rect 150102 186618 185546 186854
rect 185782 186618 185866 186854
rect 186102 186618 221546 186854
rect 221782 186618 221866 186854
rect 222102 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 588810 186854
rect -4886 186586 588810 186618
rect -2966 183454 586890 183486
rect -2966 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 244250 183454
rect 244486 183218 274970 183454
rect 275206 183218 305690 183454
rect 305926 183218 336410 183454
rect 336646 183218 367130 183454
rect 367366 183218 397850 183454
rect 398086 183218 428570 183454
rect 428806 183218 459290 183454
rect 459526 183218 490010 183454
rect 490246 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 586890 183454
rect -2966 183134 586890 183218
rect -2966 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 244250 183134
rect 244486 182898 274970 183134
rect 275206 182898 305690 183134
rect 305926 182898 336410 183134
rect 336646 182898 367130 183134
rect 367366 182898 397850 183134
rect 398086 182898 428570 183134
rect 428806 182898 459290 183134
rect 459526 182898 490010 183134
rect 490246 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 586890 183134
rect -2966 182866 586890 182898
rect -8726 176614 592650 176646
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 66986 176614
rect 67222 176378 67306 176614
rect 67542 176378 102986 176614
rect 103222 176378 103306 176614
rect 103542 176378 138986 176614
rect 139222 176378 139306 176614
rect 139542 176378 174986 176614
rect 175222 176378 175306 176614
rect 175542 176378 210986 176614
rect 211222 176378 211306 176614
rect 211542 176378 246986 176614
rect 247222 176378 247306 176614
rect 247542 176378 282986 176614
rect 283222 176378 283306 176614
rect 283542 176378 318986 176614
rect 319222 176378 319306 176614
rect 319542 176378 354986 176614
rect 355222 176378 355306 176614
rect 355542 176378 390986 176614
rect 391222 176378 391306 176614
rect 391542 176378 426986 176614
rect 427222 176378 427306 176614
rect 427542 176378 462986 176614
rect 463222 176378 463306 176614
rect 463542 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect -8726 176294 592650 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 66986 176294
rect 67222 176058 67306 176294
rect 67542 176058 102986 176294
rect 103222 176058 103306 176294
rect 103542 176058 138986 176294
rect 139222 176058 139306 176294
rect 139542 176058 174986 176294
rect 175222 176058 175306 176294
rect 175542 176058 210986 176294
rect 211222 176058 211306 176294
rect 211542 176058 246986 176294
rect 247222 176058 247306 176294
rect 247542 176058 282986 176294
rect 283222 176058 283306 176294
rect 283542 176058 318986 176294
rect 319222 176058 319306 176294
rect 319542 176058 354986 176294
rect 355222 176058 355306 176294
rect 355542 176058 390986 176294
rect 391222 176058 391306 176294
rect 391542 176058 426986 176294
rect 427222 176058 427306 176294
rect 427542 176058 462986 176294
rect 463222 176058 463306 176294
rect 463542 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect -8726 176026 592650 176058
rect -6806 172894 590730 172926
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 63266 172894
rect 63502 172658 63586 172894
rect 63822 172658 99266 172894
rect 99502 172658 99586 172894
rect 99822 172658 135266 172894
rect 135502 172658 135586 172894
rect 135822 172658 171266 172894
rect 171502 172658 171586 172894
rect 171822 172658 207266 172894
rect 207502 172658 207586 172894
rect 207822 172658 243266 172894
rect 243502 172658 243586 172894
rect 243822 172658 279266 172894
rect 279502 172658 279586 172894
rect 279822 172658 315266 172894
rect 315502 172658 315586 172894
rect 315822 172658 351266 172894
rect 351502 172658 351586 172894
rect 351822 172658 387266 172894
rect 387502 172658 387586 172894
rect 387822 172658 423266 172894
rect 423502 172658 423586 172894
rect 423822 172658 459266 172894
rect 459502 172658 459586 172894
rect 459822 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect -6806 172574 590730 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 63266 172574
rect 63502 172338 63586 172574
rect 63822 172338 99266 172574
rect 99502 172338 99586 172574
rect 99822 172338 135266 172574
rect 135502 172338 135586 172574
rect 135822 172338 171266 172574
rect 171502 172338 171586 172574
rect 171822 172338 207266 172574
rect 207502 172338 207586 172574
rect 207822 172338 243266 172574
rect 243502 172338 243586 172574
rect 243822 172338 279266 172574
rect 279502 172338 279586 172574
rect 279822 172338 315266 172574
rect 315502 172338 315586 172574
rect 315822 172338 351266 172574
rect 351502 172338 351586 172574
rect 351822 172338 387266 172574
rect 387502 172338 387586 172574
rect 387822 172338 423266 172574
rect 423502 172338 423586 172574
rect 423822 172338 459266 172574
rect 459502 172338 459586 172574
rect 459822 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect -6806 172306 590730 172338
rect -4886 169174 588810 169206
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 59546 169174
rect 59782 168938 59866 169174
rect 60102 168938 95546 169174
rect 95782 168938 95866 169174
rect 96102 168938 131546 169174
rect 131782 168938 131866 169174
rect 132102 168938 167546 169174
rect 167782 168938 167866 169174
rect 168102 168938 203546 169174
rect 203782 168938 203866 169174
rect 204102 168938 239546 169174
rect 239782 168938 239866 169174
rect 240102 168938 275546 169174
rect 275782 168938 275866 169174
rect 276102 168938 311546 169174
rect 311782 168938 311866 169174
rect 312102 168938 347546 169174
rect 347782 168938 347866 169174
rect 348102 168938 383546 169174
rect 383782 168938 383866 169174
rect 384102 168938 419546 169174
rect 419782 168938 419866 169174
rect 420102 168938 455546 169174
rect 455782 168938 455866 169174
rect 456102 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect -4886 168854 588810 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 59546 168854
rect 59782 168618 59866 168854
rect 60102 168618 95546 168854
rect 95782 168618 95866 168854
rect 96102 168618 131546 168854
rect 131782 168618 131866 168854
rect 132102 168618 167546 168854
rect 167782 168618 167866 168854
rect 168102 168618 203546 168854
rect 203782 168618 203866 168854
rect 204102 168618 239546 168854
rect 239782 168618 239866 168854
rect 240102 168618 275546 168854
rect 275782 168618 275866 168854
rect 276102 168618 311546 168854
rect 311782 168618 311866 168854
rect 312102 168618 347546 168854
rect 347782 168618 347866 168854
rect 348102 168618 383546 168854
rect 383782 168618 383866 168854
rect 384102 168618 419546 168854
rect 419782 168618 419866 168854
rect 420102 168618 455546 168854
rect 455782 168618 455866 168854
rect 456102 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect -4886 168586 588810 168618
rect -2966 165454 586890 165486
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 163826 165454
rect 164062 165218 164146 165454
rect 164382 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect -2966 165134 586890 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 163826 165134
rect 164062 164898 164146 165134
rect 164382 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect -2966 164866 586890 164898
rect -8726 158614 592650 158646
rect -8726 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 84986 158614
rect 85222 158378 85306 158614
rect 85542 158378 120986 158614
rect 121222 158378 121306 158614
rect 121542 158378 156986 158614
rect 157222 158378 157306 158614
rect 157542 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 228986 158614
rect 229222 158378 229306 158614
rect 229542 158378 264986 158614
rect 265222 158378 265306 158614
rect 265542 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 84986 158294
rect 85222 158058 85306 158294
rect 85542 158058 120986 158294
rect 121222 158058 121306 158294
rect 121542 158058 156986 158294
rect 157222 158058 157306 158294
rect 157542 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 228986 158294
rect 229222 158058 229306 158294
rect 229542 158058 264986 158294
rect 265222 158058 265306 158294
rect 265542 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 592650 158294
rect -8726 158026 592650 158058
rect -6806 154894 590730 154926
rect -6806 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 81266 154894
rect 81502 154658 81586 154894
rect 81822 154658 117266 154894
rect 117502 154658 117586 154894
rect 117822 154658 153266 154894
rect 153502 154658 153586 154894
rect 153822 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 225266 154894
rect 225502 154658 225586 154894
rect 225822 154658 261266 154894
rect 261502 154658 261586 154894
rect 261822 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 590730 154894
rect -6806 154574 590730 154658
rect -6806 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 81266 154574
rect 81502 154338 81586 154574
rect 81822 154338 117266 154574
rect 117502 154338 117586 154574
rect 117822 154338 153266 154574
rect 153502 154338 153586 154574
rect 153822 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 225266 154574
rect 225502 154338 225586 154574
rect 225822 154338 261266 154574
rect 261502 154338 261586 154574
rect 261822 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 590730 154574
rect -6806 154306 590730 154338
rect -4886 151174 588810 151206
rect -4886 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 77546 151174
rect 77782 150938 77866 151174
rect 78102 150938 113546 151174
rect 113782 150938 113866 151174
rect 114102 150938 149546 151174
rect 149782 150938 149866 151174
rect 150102 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 221546 151174
rect 221782 150938 221866 151174
rect 222102 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 588810 151174
rect -4886 150854 588810 150938
rect -4886 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 77546 150854
rect 77782 150618 77866 150854
rect 78102 150618 113546 150854
rect 113782 150618 113866 150854
rect 114102 150618 149546 150854
rect 149782 150618 149866 150854
rect 150102 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 221546 150854
rect 221782 150618 221866 150854
rect 222102 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 588810 150854
rect -4886 150586 588810 150618
rect -2966 147454 586890 147486
rect -2966 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 586890 147454
rect -2966 147134 586890 147218
rect -2966 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 586890 147134
rect -2966 146866 586890 146898
rect -8726 140614 592650 140646
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 66986 140614
rect 67222 140378 67306 140614
rect 67542 140378 102986 140614
rect 103222 140378 103306 140614
rect 103542 140378 138986 140614
rect 139222 140378 139306 140614
rect 139542 140378 174986 140614
rect 175222 140378 175306 140614
rect 175542 140378 210986 140614
rect 211222 140378 211306 140614
rect 211542 140378 246986 140614
rect 247222 140378 247306 140614
rect 247542 140378 282986 140614
rect 283222 140378 283306 140614
rect 283542 140378 318986 140614
rect 319222 140378 319306 140614
rect 319542 140378 354986 140614
rect 355222 140378 355306 140614
rect 355542 140378 390986 140614
rect 391222 140378 391306 140614
rect 391542 140378 426986 140614
rect 427222 140378 427306 140614
rect 427542 140378 462986 140614
rect 463222 140378 463306 140614
rect 463542 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect -8726 140294 592650 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 66986 140294
rect 67222 140058 67306 140294
rect 67542 140058 102986 140294
rect 103222 140058 103306 140294
rect 103542 140058 138986 140294
rect 139222 140058 139306 140294
rect 139542 140058 174986 140294
rect 175222 140058 175306 140294
rect 175542 140058 210986 140294
rect 211222 140058 211306 140294
rect 211542 140058 246986 140294
rect 247222 140058 247306 140294
rect 247542 140058 282986 140294
rect 283222 140058 283306 140294
rect 283542 140058 318986 140294
rect 319222 140058 319306 140294
rect 319542 140058 354986 140294
rect 355222 140058 355306 140294
rect 355542 140058 390986 140294
rect 391222 140058 391306 140294
rect 391542 140058 426986 140294
rect 427222 140058 427306 140294
rect 427542 140058 462986 140294
rect 463222 140058 463306 140294
rect 463542 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect -8726 140026 592650 140058
rect -6806 136894 590730 136926
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 99266 136894
rect 99502 136658 99586 136894
rect 99822 136658 135266 136894
rect 135502 136658 135586 136894
rect 135822 136658 171266 136894
rect 171502 136658 171586 136894
rect 171822 136658 207266 136894
rect 207502 136658 207586 136894
rect 207822 136658 243266 136894
rect 243502 136658 243586 136894
rect 243822 136658 279266 136894
rect 279502 136658 279586 136894
rect 279822 136658 315266 136894
rect 315502 136658 315586 136894
rect 315822 136658 351266 136894
rect 351502 136658 351586 136894
rect 351822 136658 387266 136894
rect 387502 136658 387586 136894
rect 387822 136658 423266 136894
rect 423502 136658 423586 136894
rect 423822 136658 459266 136894
rect 459502 136658 459586 136894
rect 459822 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect -6806 136574 590730 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 99266 136574
rect 99502 136338 99586 136574
rect 99822 136338 135266 136574
rect 135502 136338 135586 136574
rect 135822 136338 171266 136574
rect 171502 136338 171586 136574
rect 171822 136338 207266 136574
rect 207502 136338 207586 136574
rect 207822 136338 243266 136574
rect 243502 136338 243586 136574
rect 243822 136338 279266 136574
rect 279502 136338 279586 136574
rect 279822 136338 315266 136574
rect 315502 136338 315586 136574
rect 315822 136338 351266 136574
rect 351502 136338 351586 136574
rect 351822 136338 387266 136574
rect 387502 136338 387586 136574
rect 387822 136338 423266 136574
rect 423502 136338 423586 136574
rect 423822 136338 459266 136574
rect 459502 136338 459586 136574
rect 459822 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect -6806 136306 590730 136338
rect -4886 133174 588810 133206
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 95546 133174
rect 95782 132938 95866 133174
rect 96102 132938 131546 133174
rect 131782 132938 131866 133174
rect 132102 132938 167546 133174
rect 167782 132938 167866 133174
rect 168102 132938 203546 133174
rect 203782 132938 203866 133174
rect 204102 132938 239546 133174
rect 239782 132938 239866 133174
rect 240102 132938 275546 133174
rect 275782 132938 275866 133174
rect 276102 132938 311546 133174
rect 311782 132938 311866 133174
rect 312102 132938 347546 133174
rect 347782 132938 347866 133174
rect 348102 132938 383546 133174
rect 383782 132938 383866 133174
rect 384102 132938 419546 133174
rect 419782 132938 419866 133174
rect 420102 132938 455546 133174
rect 455782 132938 455866 133174
rect 456102 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect -4886 132854 588810 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 95546 132854
rect 95782 132618 95866 132854
rect 96102 132618 131546 132854
rect 131782 132618 131866 132854
rect 132102 132618 167546 132854
rect 167782 132618 167866 132854
rect 168102 132618 203546 132854
rect 203782 132618 203866 132854
rect 204102 132618 239546 132854
rect 239782 132618 239866 132854
rect 240102 132618 275546 132854
rect 275782 132618 275866 132854
rect 276102 132618 311546 132854
rect 311782 132618 311866 132854
rect 312102 132618 347546 132854
rect 347782 132618 347866 132854
rect 348102 132618 383546 132854
rect 383782 132618 383866 132854
rect 384102 132618 419546 132854
rect 419782 132618 419866 132854
rect 420102 132618 455546 132854
rect 455782 132618 455866 132854
rect 456102 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect -4886 132586 588810 132618
rect -2966 129454 586890 129486
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 127826 129454
rect 128062 129218 128146 129454
rect 128382 129218 163826 129454
rect 164062 129218 164146 129454
rect 164382 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect -2966 129134 586890 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 127826 129134
rect 128062 128898 128146 129134
rect 128382 128898 163826 129134
rect 164062 128898 164146 129134
rect 164382 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect -2966 128866 586890 128898
rect -8726 122614 592650 122646
rect -8726 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 84986 122614
rect 85222 122378 85306 122614
rect 85542 122378 120986 122614
rect 121222 122378 121306 122614
rect 121542 122378 156986 122614
rect 157222 122378 157306 122614
rect 157542 122378 192986 122614
rect 193222 122378 193306 122614
rect 193542 122378 228986 122614
rect 229222 122378 229306 122614
rect 229542 122378 264986 122614
rect 265222 122378 265306 122614
rect 265542 122378 300986 122614
rect 301222 122378 301306 122614
rect 301542 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 84986 122294
rect 85222 122058 85306 122294
rect 85542 122058 120986 122294
rect 121222 122058 121306 122294
rect 121542 122058 156986 122294
rect 157222 122058 157306 122294
rect 157542 122058 192986 122294
rect 193222 122058 193306 122294
rect 193542 122058 228986 122294
rect 229222 122058 229306 122294
rect 229542 122058 264986 122294
rect 265222 122058 265306 122294
rect 265542 122058 300986 122294
rect 301222 122058 301306 122294
rect 301542 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 592650 122294
rect -8726 122026 592650 122058
rect -6806 118894 590730 118926
rect -6806 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 81266 118894
rect 81502 118658 81586 118894
rect 81822 118658 117266 118894
rect 117502 118658 117586 118894
rect 117822 118658 153266 118894
rect 153502 118658 153586 118894
rect 153822 118658 189266 118894
rect 189502 118658 189586 118894
rect 189822 118658 225266 118894
rect 225502 118658 225586 118894
rect 225822 118658 261266 118894
rect 261502 118658 261586 118894
rect 261822 118658 297266 118894
rect 297502 118658 297586 118894
rect 297822 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 590730 118894
rect -6806 118574 590730 118658
rect -6806 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 81266 118574
rect 81502 118338 81586 118574
rect 81822 118338 117266 118574
rect 117502 118338 117586 118574
rect 117822 118338 153266 118574
rect 153502 118338 153586 118574
rect 153822 118338 189266 118574
rect 189502 118338 189586 118574
rect 189822 118338 225266 118574
rect 225502 118338 225586 118574
rect 225822 118338 261266 118574
rect 261502 118338 261586 118574
rect 261822 118338 297266 118574
rect 297502 118338 297586 118574
rect 297822 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 590730 118574
rect -6806 118306 590730 118338
rect -4886 115174 588810 115206
rect -4886 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 77546 115174
rect 77782 114938 77866 115174
rect 78102 114938 113546 115174
rect 113782 114938 113866 115174
rect 114102 114938 149546 115174
rect 149782 114938 149866 115174
rect 150102 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 221546 115174
rect 221782 114938 221866 115174
rect 222102 114938 257546 115174
rect 257782 114938 257866 115174
rect 258102 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 588810 115174
rect -4886 114854 588810 114938
rect -4886 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 77546 114854
rect 77782 114618 77866 114854
rect 78102 114618 113546 114854
rect 113782 114618 113866 114854
rect 114102 114618 149546 114854
rect 149782 114618 149866 114854
rect 150102 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 221546 114854
rect 221782 114618 221866 114854
rect 222102 114618 257546 114854
rect 257782 114618 257866 114854
rect 258102 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 588810 114854
rect -4886 114586 588810 114618
rect -2966 111454 586890 111486
rect -2966 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 586890 111454
rect -2966 111134 586890 111218
rect -2966 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 586890 111134
rect -2966 110866 586890 110898
rect -8726 104614 592650 104646
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 66986 104614
rect 67222 104378 67306 104614
rect 67542 104378 102986 104614
rect 103222 104378 103306 104614
rect 103542 104378 138986 104614
rect 139222 104378 139306 104614
rect 139542 104378 174986 104614
rect 175222 104378 175306 104614
rect 175542 104378 210986 104614
rect 211222 104378 211306 104614
rect 211542 104378 246986 104614
rect 247222 104378 247306 104614
rect 247542 104378 282986 104614
rect 283222 104378 283306 104614
rect 283542 104378 318986 104614
rect 319222 104378 319306 104614
rect 319542 104378 354986 104614
rect 355222 104378 355306 104614
rect 355542 104378 390986 104614
rect 391222 104378 391306 104614
rect 391542 104378 426986 104614
rect 427222 104378 427306 104614
rect 427542 104378 462986 104614
rect 463222 104378 463306 104614
rect 463542 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect -8726 104294 592650 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 66986 104294
rect 67222 104058 67306 104294
rect 67542 104058 102986 104294
rect 103222 104058 103306 104294
rect 103542 104058 138986 104294
rect 139222 104058 139306 104294
rect 139542 104058 174986 104294
rect 175222 104058 175306 104294
rect 175542 104058 210986 104294
rect 211222 104058 211306 104294
rect 211542 104058 246986 104294
rect 247222 104058 247306 104294
rect 247542 104058 282986 104294
rect 283222 104058 283306 104294
rect 283542 104058 318986 104294
rect 319222 104058 319306 104294
rect 319542 104058 354986 104294
rect 355222 104058 355306 104294
rect 355542 104058 390986 104294
rect 391222 104058 391306 104294
rect 391542 104058 426986 104294
rect 427222 104058 427306 104294
rect 427542 104058 462986 104294
rect 463222 104058 463306 104294
rect 463542 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect -8726 104026 592650 104058
rect -6806 100894 590730 100926
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 63266 100894
rect 63502 100658 63586 100894
rect 63822 100658 99266 100894
rect 99502 100658 99586 100894
rect 99822 100658 135266 100894
rect 135502 100658 135586 100894
rect 135822 100658 171266 100894
rect 171502 100658 171586 100894
rect 171822 100658 207266 100894
rect 207502 100658 207586 100894
rect 207822 100658 243266 100894
rect 243502 100658 243586 100894
rect 243822 100658 279266 100894
rect 279502 100658 279586 100894
rect 279822 100658 315266 100894
rect 315502 100658 315586 100894
rect 315822 100658 351266 100894
rect 351502 100658 351586 100894
rect 351822 100658 387266 100894
rect 387502 100658 387586 100894
rect 387822 100658 423266 100894
rect 423502 100658 423586 100894
rect 423822 100658 459266 100894
rect 459502 100658 459586 100894
rect 459822 100658 495266 100894
rect 495502 100658 495586 100894
rect 495822 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect -6806 100574 590730 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 63266 100574
rect 63502 100338 63586 100574
rect 63822 100338 99266 100574
rect 99502 100338 99586 100574
rect 99822 100338 135266 100574
rect 135502 100338 135586 100574
rect 135822 100338 171266 100574
rect 171502 100338 171586 100574
rect 171822 100338 207266 100574
rect 207502 100338 207586 100574
rect 207822 100338 243266 100574
rect 243502 100338 243586 100574
rect 243822 100338 279266 100574
rect 279502 100338 279586 100574
rect 279822 100338 315266 100574
rect 315502 100338 315586 100574
rect 315822 100338 351266 100574
rect 351502 100338 351586 100574
rect 351822 100338 387266 100574
rect 387502 100338 387586 100574
rect 387822 100338 423266 100574
rect 423502 100338 423586 100574
rect 423822 100338 459266 100574
rect 459502 100338 459586 100574
rect 459822 100338 495266 100574
rect 495502 100338 495586 100574
rect 495822 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect -6806 100306 590730 100338
rect -4886 97174 588810 97206
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 59546 97174
rect 59782 96938 59866 97174
rect 60102 96938 95546 97174
rect 95782 96938 95866 97174
rect 96102 96938 131546 97174
rect 131782 96938 131866 97174
rect 132102 96938 167546 97174
rect 167782 96938 167866 97174
rect 168102 96938 203546 97174
rect 203782 96938 203866 97174
rect 204102 96938 239546 97174
rect 239782 96938 239866 97174
rect 240102 96938 275546 97174
rect 275782 96938 275866 97174
rect 276102 96938 311546 97174
rect 311782 96938 311866 97174
rect 312102 96938 347546 97174
rect 347782 96938 347866 97174
rect 348102 96938 383546 97174
rect 383782 96938 383866 97174
rect 384102 96938 419546 97174
rect 419782 96938 419866 97174
rect 420102 96938 455546 97174
rect 455782 96938 455866 97174
rect 456102 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect -4886 96854 588810 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 59546 96854
rect 59782 96618 59866 96854
rect 60102 96618 95546 96854
rect 95782 96618 95866 96854
rect 96102 96618 131546 96854
rect 131782 96618 131866 96854
rect 132102 96618 167546 96854
rect 167782 96618 167866 96854
rect 168102 96618 203546 96854
rect 203782 96618 203866 96854
rect 204102 96618 239546 96854
rect 239782 96618 239866 96854
rect 240102 96618 275546 96854
rect 275782 96618 275866 96854
rect 276102 96618 311546 96854
rect 311782 96618 311866 96854
rect 312102 96618 347546 96854
rect 347782 96618 347866 96854
rect 348102 96618 383546 96854
rect 383782 96618 383866 96854
rect 384102 96618 419546 96854
rect 419782 96618 419866 96854
rect 420102 96618 455546 96854
rect 455782 96618 455866 96854
rect 456102 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect -4886 96586 588810 96618
rect -2966 93454 586890 93486
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 127826 93454
rect 128062 93218 128146 93454
rect 128382 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect -2966 93134 586890 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 127826 93134
rect 128062 92898 128146 93134
rect 128382 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect -2966 92866 586890 92898
rect -8726 86614 592650 86646
rect -8726 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 120986 86614
rect 121222 86378 121306 86614
rect 121542 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 192986 86614
rect 193222 86378 193306 86614
rect 193542 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 120986 86294
rect 121222 86058 121306 86294
rect 121542 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 192986 86294
rect 193222 86058 193306 86294
rect 193542 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 592650 86294
rect -8726 86026 592650 86058
rect -6806 82894 590730 82926
rect -6806 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 117266 82894
rect 117502 82658 117586 82894
rect 117822 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 189266 82894
rect 189502 82658 189586 82894
rect 189822 82658 225266 82894
rect 225502 82658 225586 82894
rect 225822 82658 261266 82894
rect 261502 82658 261586 82894
rect 261822 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 590730 82894
rect -6806 82574 590730 82658
rect -6806 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 117266 82574
rect 117502 82338 117586 82574
rect 117822 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 189266 82574
rect 189502 82338 189586 82574
rect 189822 82338 225266 82574
rect 225502 82338 225586 82574
rect 225822 82338 261266 82574
rect 261502 82338 261586 82574
rect 261822 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 590730 82574
rect -6806 82306 590730 82338
rect -4886 79174 588810 79206
rect -4886 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 588810 79174
rect -4886 78854 588810 78938
rect -4886 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 588810 78854
rect -4886 78586 588810 78618
rect -2966 75454 586890 75486
rect -2966 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 586890 75454
rect -2966 75134 586890 75218
rect -2966 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 586890 75134
rect -2966 74866 586890 74898
rect -8726 68614 592650 68646
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 66986 68614
rect 67222 68378 67306 68614
rect 67542 68378 102986 68614
rect 103222 68378 103306 68614
rect 103542 68378 138986 68614
rect 139222 68378 139306 68614
rect 139542 68378 174986 68614
rect 175222 68378 175306 68614
rect 175542 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 246986 68614
rect 247222 68378 247306 68614
rect 247542 68378 282986 68614
rect 283222 68378 283306 68614
rect 283542 68378 318986 68614
rect 319222 68378 319306 68614
rect 319542 68378 354986 68614
rect 355222 68378 355306 68614
rect 355542 68378 390986 68614
rect 391222 68378 391306 68614
rect 391542 68378 426986 68614
rect 427222 68378 427306 68614
rect 427542 68378 462986 68614
rect 463222 68378 463306 68614
rect 463542 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect -8726 68294 592650 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 66986 68294
rect 67222 68058 67306 68294
rect 67542 68058 102986 68294
rect 103222 68058 103306 68294
rect 103542 68058 138986 68294
rect 139222 68058 139306 68294
rect 139542 68058 174986 68294
rect 175222 68058 175306 68294
rect 175542 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 246986 68294
rect 247222 68058 247306 68294
rect 247542 68058 282986 68294
rect 283222 68058 283306 68294
rect 283542 68058 318986 68294
rect 319222 68058 319306 68294
rect 319542 68058 354986 68294
rect 355222 68058 355306 68294
rect 355542 68058 390986 68294
rect 391222 68058 391306 68294
rect 391542 68058 426986 68294
rect 427222 68058 427306 68294
rect 427542 68058 462986 68294
rect 463222 68058 463306 68294
rect 463542 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect -8726 68026 592650 68058
rect -6806 64894 590730 64926
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 63266 64894
rect 63502 64658 63586 64894
rect 63822 64658 99266 64894
rect 99502 64658 99586 64894
rect 99822 64658 135266 64894
rect 135502 64658 135586 64894
rect 135822 64658 171266 64894
rect 171502 64658 171586 64894
rect 171822 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 243266 64894
rect 243502 64658 243586 64894
rect 243822 64658 279266 64894
rect 279502 64658 279586 64894
rect 279822 64658 315266 64894
rect 315502 64658 315586 64894
rect 315822 64658 351266 64894
rect 351502 64658 351586 64894
rect 351822 64658 387266 64894
rect 387502 64658 387586 64894
rect 387822 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect -6806 64574 590730 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 63266 64574
rect 63502 64338 63586 64574
rect 63822 64338 99266 64574
rect 99502 64338 99586 64574
rect 99822 64338 135266 64574
rect 135502 64338 135586 64574
rect 135822 64338 171266 64574
rect 171502 64338 171586 64574
rect 171822 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 243266 64574
rect 243502 64338 243586 64574
rect 243822 64338 279266 64574
rect 279502 64338 279586 64574
rect 279822 64338 315266 64574
rect 315502 64338 315586 64574
rect 315822 64338 351266 64574
rect 351502 64338 351586 64574
rect 351822 64338 387266 64574
rect 387502 64338 387586 64574
rect 387822 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect -6806 64306 590730 64338
rect -4886 61174 588810 61206
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 59546 61174
rect 59782 60938 59866 61174
rect 60102 60938 95546 61174
rect 95782 60938 95866 61174
rect 96102 60938 131546 61174
rect 131782 60938 131866 61174
rect 132102 60938 167546 61174
rect 167782 60938 167866 61174
rect 168102 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 239546 61174
rect 239782 60938 239866 61174
rect 240102 60938 275546 61174
rect 275782 60938 275866 61174
rect 276102 60938 311546 61174
rect 311782 60938 311866 61174
rect 312102 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect -4886 60854 588810 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 59546 60854
rect 59782 60618 59866 60854
rect 60102 60618 95546 60854
rect 95782 60618 95866 60854
rect 96102 60618 131546 60854
rect 131782 60618 131866 60854
rect 132102 60618 167546 60854
rect 167782 60618 167866 60854
rect 168102 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 239546 60854
rect 239782 60618 239866 60854
rect 240102 60618 275546 60854
rect 275782 60618 275866 60854
rect 276102 60618 311546 60854
rect 311782 60618 311866 60854
rect 312102 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect -4886 60586 588810 60618
rect -2966 57454 586890 57486
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect -2966 57134 586890 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect -2966 56866 586890 56898
rect -8726 50614 592650 50646
rect -8726 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 592650 50294
rect -8726 50026 592650 50058
rect -6806 46894 590730 46926
rect -6806 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 590730 46894
rect -6806 46574 590730 46658
rect -6806 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 590730 46574
rect -6806 46306 590730 46338
rect -4886 43174 588810 43206
rect -4886 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 588810 43174
rect -4886 42854 588810 42938
rect -4886 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 588810 42854
rect -4886 42586 588810 42618
rect -2966 39454 586890 39486
rect -2966 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 586890 39454
rect -2966 39134 586890 39218
rect -2966 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 586890 39134
rect -2966 38866 586890 38898
rect -8726 32614 592650 32646
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect -8726 32294 592650 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect -8726 32026 592650 32058
rect -6806 28894 590730 28926
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect -6806 28574 590730 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect -6806 28306 590730 28338
rect -4886 25174 588810 25206
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect -4886 24854 588810 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect -4886 24586 588810 24618
rect -2966 21454 586890 21486
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect -2966 21134 586890 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect -2966 20866 586890 20898
rect -8726 14614 592650 14646
rect -8726 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 592650 14294
rect -8726 14026 592650 14058
rect -6806 10894 590730 10926
rect -6806 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 590730 10894
rect -6806 10574 590730 10658
rect -6806 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 590730 10574
rect -6806 10306 590730 10338
rect -4886 7174 588810 7206
rect -4886 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 588810 7174
rect -4886 6854 588810 6938
rect -4886 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 588810 6854
rect -4886 6586 588810 6618
rect -2966 3454 586890 3486
rect -2966 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 586890 3454
rect -2966 3134 586890 3218
rect -2966 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 586890 3134
rect -2966 2866 586890 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use sky130_sram_2kbyte_1rw1r_32x512_8  BB_SRAM
timestamp 0
transform 1 0 50000 0 1 380000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  VB_SRAM
timestamp 0
transform 1 0 50000 0 1 200000
box 0 0 136620 83308
use c0_system  mprj
timestamp 0
transform 1 0 240000 0 1 180000
box 0 0 258888 259616
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 38866 586890 39486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 74866 586890 75486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 110866 586890 111486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 146866 586890 147486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 182866 586890 183486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 218866 586890 219486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 254866 586890 255486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 290866 586890 291486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 326866 586890 327486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 362866 586890 363486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 398866 586890 399486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 434866 586890 435486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 470866 586890 471486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 578866 586890 579486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 614866 586890 615486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 650866 586890 651486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 686866 586890 687486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 -1894 254414 178000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 -1894 290414 178000 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 -1894 326414 178000 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 -1894 362414 178000 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 -1894 398414 178000 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 -1894 434414 178000 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 -1894 470414 178000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 -1894 74414 198000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 -1894 110414 198000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 -1894 146414 198000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 -1894 182414 198000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 285308 74414 378000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 285308 110414 378000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 285308 146414 378000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 285308 182414 378000 6 vccd1
port 531 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 1794 -1894 2414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 -1894 38414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 465308 74414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 465308 110414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 465308 146414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 465308 182414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 -1894 218414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 442000 254414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 442000 290414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 442000 326414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 442000 362414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 442000 398414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 442000 434414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 442000 470414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 -1894 506414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 -1894 542414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 577794 -1894 578414 705830 6 vccd1
port 531 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 532 nsew power input
rlabel metal5 s -4886 6586 588810 7206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 42586 588810 43206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 78586 588810 79206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 114586 588810 115206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 150586 588810 151206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 186586 588810 187206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 222586 588810 223206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 258586 588810 259206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 294586 588810 295206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 330586 588810 331206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 366586 588810 367206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 402586 588810 403206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 438586 588810 439206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 474586 588810 475206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 510586 588810 511206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 546586 588810 547206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 582586 588810 583206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 618586 588810 619206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 654586 588810 655206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 690586 588810 691206 6 vccd2
port 532 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 -3814 258134 178000 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 -3814 294134 178000 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 -3814 330134 178000 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 -3814 366134 178000 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 -3814 402134 178000 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 -3814 438134 178000 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 -3814 474134 178000 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 -3814 78134 198000 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 -3814 114134 198000 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 -3814 150134 198000 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 -3814 186134 198000 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 285308 78134 378000 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 285308 114134 378000 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 285308 150134 378000 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 285308 186134 378000 6 vccd2
port 532 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 532 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 5514 -3814 6134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 41514 -3814 42134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 465308 78134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 465308 114134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 465308 150134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 465308 186134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 -3814 222134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 442000 258134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 442000 294134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 442000 330134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 442000 366134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 442000 402134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 442000 438134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 442000 474134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 -3814 510134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 545514 -3814 546134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 581514 -3814 582134 707750 6 vccd2
port 532 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 533 nsew power input
rlabel metal5 s -6806 10306 590730 10926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 46306 590730 46926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 82306 590730 82926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 118306 590730 118926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 154306 590730 154926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 190306 590730 190926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 226306 590730 226926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 262306 590730 262926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 298306 590730 298926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 334306 590730 334926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 370306 590730 370926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 406306 590730 406926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 442306 590730 442926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 478306 590730 478926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 514306 590730 514926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 550306 590730 550926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 586306 590730 586926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 622306 590730 622926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 658306 590730 658926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 694306 590730 694926 6 vdda1
port 533 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 -5734 261854 178000 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 -5734 297854 178000 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 -5734 333854 178000 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 -5734 369854 178000 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 -5734 405854 178000 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 -5734 441854 178000 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 -5734 477854 178000 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 -5734 81854 198000 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 -5734 117854 198000 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 -5734 153854 198000 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 285308 81854 378000 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 285308 117854 378000 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 285308 153854 378000 6 vdda1
port 533 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 533 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 9234 -5734 9854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 45234 -5734 45854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 465308 81854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 465308 117854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 465308 153854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 -5734 189854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 -5734 225854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 442000 261854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 442000 297854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 442000 333854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 442000 369854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 442000 405854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 442000 441854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 442000 477854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 -5734 513854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 549234 -5734 549854 709670 6 vdda1
port 533 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 534 nsew power input
rlabel metal5 s -8726 14026 592650 14646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 50026 592650 50646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 86026 592650 86646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 122026 592650 122646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 158026 592650 158646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 194026 592650 194646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 230026 592650 230646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 266026 592650 266646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 302026 592650 302646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 338026 592650 338646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 374026 592650 374646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 410026 592650 410646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 446026 592650 446646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 482026 592650 482646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 518026 592650 518646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 554026 592650 554646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 590026 592650 590646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 626026 592650 626646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 662026 592650 662646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 698026 592650 698646 6 vdda2
port 534 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 -7654 265574 178000 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 -7654 301574 178000 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 -7654 337574 178000 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 -7654 373574 178000 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 -7654 409574 178000 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 -7654 445574 178000 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 -7654 481574 178000 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 -7654 49574 198000 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 -7654 85574 198000 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 -7654 121574 198000 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 -7654 157574 198000 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 285308 49574 378000 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 285308 85574 378000 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 285308 121574 378000 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 285308 157574 378000 6 vdda2
port 534 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 534 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 12954 -7654 13574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 465308 49574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 465308 85574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 465308 121574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 465308 157574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 -7654 193574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 -7654 229574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 442000 265574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 442000 301574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 442000 337574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 442000 373574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 442000 409574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 442000 445574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 442000 481574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 -7654 517574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 552954 -7654 553574 711590 6 vdda2
port 534 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 28306 590730 28926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 64306 590730 64926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 100306 590730 100926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 136306 590730 136926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 172306 590730 172926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 208306 590730 208926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 244306 590730 244926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 280306 590730 280926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 316306 590730 316926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 352306 590730 352926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 388306 590730 388926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 424306 590730 424926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 460306 590730 460926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 496306 590730 496926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 532306 590730 532926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 568306 590730 568926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 604306 590730 604926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 640306 590730 640926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 676306 590730 676926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 -5734 243854 178000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 -5734 279854 178000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 -5734 315854 178000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 -5734 351854 178000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 -5734 387854 178000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 -5734 423854 178000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 -5734 459854 178000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 -5734 495854 178000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 -5734 63854 198000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 -5734 99854 198000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 -5734 135854 198000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 -5734 171854 198000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 285308 63854 378000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 285308 99854 378000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 285308 135854 378000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 285308 171854 378000 6 vssa1
port 535 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 535 nsew ground input
rlabel metal4 s 27234 -5734 27854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 465308 63854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 465308 99854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 465308 135854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 465308 171854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 -5734 207854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 442000 243854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 442000 279854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 442000 315854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 442000 351854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 442000 387854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 442000 423854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 442000 459854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 442000 495854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 -5734 531854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 567234 -5734 567854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 32026 592650 32646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 68026 592650 68646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 104026 592650 104646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 140026 592650 140646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 176026 592650 176646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 212026 592650 212646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 248026 592650 248646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 284026 592650 284646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 320026 592650 320646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 356026 592650 356646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 392026 592650 392646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 428026 592650 428646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 464026 592650 464646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 500026 592650 500646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 536026 592650 536646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 572026 592650 572646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 608026 592650 608646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 644026 592650 644646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 680026 592650 680646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 -7654 247574 178000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 -7654 283574 178000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 -7654 319574 178000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 -7654 355574 178000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 -7654 391574 178000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 -7654 427574 178000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 -7654 463574 178000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 -7654 499574 178000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 -7654 67574 198000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 -7654 103574 198000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 -7654 139574 198000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 -7654 175574 198000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 285308 67574 378000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 285308 103574 378000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 285308 139574 378000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 285308 175574 378000 6 vssa2
port 536 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 -7654 31574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 465308 67574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 465308 103574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 465308 139574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 465308 175574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 -7654 211574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 442000 247574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 442000 283574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 442000 319574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 442000 355574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 442000 391574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 442000 427574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 442000 463574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 442000 499574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 -7654 535574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 570954 -7654 571574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 20866 586890 21486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 56866 586890 57486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 92866 586890 93486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 128866 586890 129486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 164866 586890 165486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 200866 586890 201486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 236866 586890 237486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 272866 586890 273486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 308866 586890 309486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 344866 586890 345486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 380866 586890 381486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 416866 586890 417486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 452866 586890 453486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 488866 586890 489486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 524866 586890 525486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 560866 586890 561486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 596866 586890 597486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 632866 586890 633486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 668866 586890 669486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 -1894 272414 178000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 -1894 308414 178000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 -1894 344414 178000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 -1894 380414 178000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 -1894 416414 178000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 -1894 452414 178000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 -1894 488414 178000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 -1894 56414 198000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 -1894 92414 198000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 -1894 128414 198000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 -1894 164414 198000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 285308 56414 378000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 285308 92414 378000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 285308 128414 378000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 285308 164414 378000 6 vssd1
port 537 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 537 nsew ground input
rlabel metal4 s 19794 -1894 20414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 465308 56414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 465308 92414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 465308 128414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 465308 164414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 -1894 200414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 -1894 236414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 442000 272414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 442000 308414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 442000 344414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 442000 380414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 442000 416414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 442000 452414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 442000 488414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 -1894 524414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 559794 -1894 560414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 24586 588810 25206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 60586 588810 61206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 96586 588810 97206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 132586 588810 133206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 168586 588810 169206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 204586 588810 205206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 240586 588810 241206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 276586 588810 277206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 312586 588810 313206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 348586 588810 349206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 384586 588810 385206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 420586 588810 421206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 456586 588810 457206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 492586 588810 493206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 528586 588810 529206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 564586 588810 565206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 600586 588810 601206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 636586 588810 637206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 672586 588810 673206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 -3814 240134 178000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 -3814 276134 178000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 -3814 312134 178000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 -3814 348134 178000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 -3814 384134 178000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 -3814 420134 178000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 -3814 456134 178000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 -3814 492134 178000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 -3814 60134 198000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 -3814 96134 198000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 -3814 132134 198000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 -3814 168134 198000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 285308 60134 378000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 285308 96134 378000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 285308 132134 378000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 285308 168134 378000 6 vssd2
port 538 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 538 nsew ground input
rlabel metal4 s 23514 -3814 24134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 465308 60134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 465308 96134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 465308 132134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 465308 168134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 -3814 204134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 442000 240134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 442000 276134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 442000 312134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 442000 348134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 442000 384134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 442000 420134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 442000 456134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 442000 492134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 -3814 528134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 563514 -3814 564134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 541 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 607 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 608 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 609 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 610 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 611 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 612 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 613 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 614 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 615 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 616 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 617 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 618 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 619 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 620 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 621 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 622 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 623 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 624 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 625 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 626 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 627 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 628 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 629 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 630 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 631 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 632 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 633 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 634 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 635 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 636 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 637 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 638 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1647715346
<< obsli1 >>
rect 1104 2159 238832 357425
<< obsm1 >>
rect 750 2128 238832 357456
<< metal2 >>
rect 1582 0 1638 800
rect 4710 0 4766 800
rect 7930 0 7986 800
rect 11150 0 11206 800
rect 14370 0 14426 800
rect 17498 0 17554 800
rect 20718 0 20774 800
rect 23938 0 23994 800
rect 27158 0 27214 800
rect 30378 0 30434 800
rect 33506 0 33562 800
rect 36726 0 36782 800
rect 39946 0 40002 800
rect 43166 0 43222 800
rect 46386 0 46442 800
rect 49514 0 49570 800
rect 52734 0 52790 800
rect 55954 0 56010 800
rect 59174 0 59230 800
rect 62302 0 62358 800
rect 65522 0 65578 800
rect 68742 0 68798 800
rect 71962 0 72018 800
rect 75182 0 75238 800
rect 78310 0 78366 800
rect 81530 0 81586 800
rect 84750 0 84806 800
rect 87970 0 88026 800
rect 91190 0 91246 800
rect 94318 0 94374 800
rect 97538 0 97594 800
rect 100758 0 100814 800
rect 103978 0 104034 800
rect 107106 0 107162 800
rect 110326 0 110382 800
rect 113546 0 113602 800
rect 116766 0 116822 800
rect 119986 0 120042 800
rect 123114 0 123170 800
rect 126334 0 126390 800
rect 129554 0 129610 800
rect 132774 0 132830 800
rect 135994 0 136050 800
rect 139122 0 139178 800
rect 142342 0 142398 800
rect 145562 0 145618 800
rect 148782 0 148838 800
rect 151910 0 151966 800
rect 155130 0 155186 800
rect 158350 0 158406 800
rect 161570 0 161626 800
rect 164790 0 164846 800
rect 167918 0 167974 800
rect 171138 0 171194 800
rect 174358 0 174414 800
rect 177578 0 177634 800
rect 180798 0 180854 800
rect 183926 0 183982 800
rect 187146 0 187202 800
rect 190366 0 190422 800
rect 193586 0 193642 800
rect 196714 0 196770 800
rect 199934 0 199990 800
rect 203154 0 203210 800
rect 206374 0 206430 800
rect 209594 0 209650 800
rect 212722 0 212778 800
rect 215942 0 215998 800
rect 219162 0 219218 800
rect 222382 0 222438 800
rect 225602 0 225658 800
rect 228730 0 228786 800
rect 231950 0 232006 800
rect 235170 0 235226 800
rect 238390 0 238446 800
<< obsm2 >>
rect 756 856 238444 359417
rect 756 575 1526 856
rect 1694 575 4654 856
rect 4822 575 7874 856
rect 8042 575 11094 856
rect 11262 575 14314 856
rect 14482 575 17442 856
rect 17610 575 20662 856
rect 20830 575 23882 856
rect 24050 575 27102 856
rect 27270 575 30322 856
rect 30490 575 33450 856
rect 33618 575 36670 856
rect 36838 575 39890 856
rect 40058 575 43110 856
rect 43278 575 46330 856
rect 46498 575 49458 856
rect 49626 575 52678 856
rect 52846 575 55898 856
rect 56066 575 59118 856
rect 59286 575 62246 856
rect 62414 575 65466 856
rect 65634 575 68686 856
rect 68854 575 71906 856
rect 72074 575 75126 856
rect 75294 575 78254 856
rect 78422 575 81474 856
rect 81642 575 84694 856
rect 84862 575 87914 856
rect 88082 575 91134 856
rect 91302 575 94262 856
rect 94430 575 97482 856
rect 97650 575 100702 856
rect 100870 575 103922 856
rect 104090 575 107050 856
rect 107218 575 110270 856
rect 110438 575 113490 856
rect 113658 575 116710 856
rect 116878 575 119930 856
rect 120098 575 123058 856
rect 123226 575 126278 856
rect 126446 575 129498 856
rect 129666 575 132718 856
rect 132886 575 135938 856
rect 136106 575 139066 856
rect 139234 575 142286 856
rect 142454 575 145506 856
rect 145674 575 148726 856
rect 148894 575 151854 856
rect 152022 575 155074 856
rect 155242 575 158294 856
rect 158462 575 161514 856
rect 161682 575 164734 856
rect 164902 575 167862 856
rect 168030 575 171082 856
rect 171250 575 174302 856
rect 174470 575 177522 856
rect 177690 575 180742 856
rect 180910 575 183870 856
rect 184038 575 187090 856
rect 187258 575 190310 856
rect 190478 575 193530 856
rect 193698 575 196658 856
rect 196826 575 199878 856
rect 200046 575 203098 856
rect 203266 575 206318 856
rect 206486 575 209538 856
rect 209706 575 212666 856
rect 212834 575 215886 856
rect 216054 575 219106 856
rect 219274 575 222326 856
rect 222494 575 225546 856
rect 225714 575 228674 856
rect 228842 575 231894 856
rect 232062 575 235114 856
rect 235282 575 238334 856
<< metal3 >>
rect 0 359320 800 359440
rect 0 358096 800 358216
rect 0 356872 800 356992
rect 0 355648 800 355768
rect 0 354424 800 354544
rect 0 353200 800 353320
rect 0 351976 800 352096
rect 0 350752 800 350872
rect 0 349528 800 349648
rect 0 348304 800 348424
rect 0 347080 800 347200
rect 0 345856 800 345976
rect 0 344632 800 344752
rect 0 343408 800 343528
rect 0 342184 800 342304
rect 0 340960 800 341080
rect 0 339736 800 339856
rect 0 338648 800 338768
rect 0 337424 800 337544
rect 0 336200 800 336320
rect 0 334976 800 335096
rect 0 333752 800 333872
rect 0 332528 800 332648
rect 0 331304 800 331424
rect 0 330080 800 330200
rect 0 328856 800 328976
rect 0 327632 800 327752
rect 0 326408 800 326528
rect 0 325184 800 325304
rect 0 323960 800 324080
rect 0 322736 800 322856
rect 0 321512 800 321632
rect 0 320288 800 320408
rect 0 319064 800 319184
rect 0 317976 800 318096
rect 0 316752 800 316872
rect 0 315528 800 315648
rect 0 314304 800 314424
rect 0 313080 800 313200
rect 0 311856 800 311976
rect 0 310632 800 310752
rect 0 309408 800 309528
rect 0 308184 800 308304
rect 0 306960 800 307080
rect 0 305736 800 305856
rect 0 304512 800 304632
rect 0 303288 800 303408
rect 0 302064 800 302184
rect 0 300840 800 300960
rect 0 299616 800 299736
rect 0 298392 800 298512
rect 0 297168 800 297288
rect 0 296080 800 296200
rect 0 294856 800 294976
rect 0 293632 800 293752
rect 0 292408 800 292528
rect 0 291184 800 291304
rect 0 289960 800 290080
rect 0 288736 800 288856
rect 0 287512 800 287632
rect 0 286288 800 286408
rect 0 285064 800 285184
rect 0 283840 800 283960
rect 0 282616 800 282736
rect 0 281392 800 281512
rect 0 280168 800 280288
rect 0 278944 800 279064
rect 0 277720 800 277840
rect 0 276496 800 276616
rect 0 275408 800 275528
rect 0 274184 800 274304
rect 0 272960 800 273080
rect 0 271736 800 271856
rect 0 270512 800 270632
rect 0 269288 800 269408
rect 0 268064 800 268184
rect 0 266840 800 266960
rect 0 265616 800 265736
rect 0 264392 800 264512
rect 0 263168 800 263288
rect 0 261944 800 262064
rect 0 260720 800 260840
rect 0 259496 800 259616
rect 0 258272 800 258392
rect 0 257048 800 257168
rect 0 255824 800 255944
rect 0 254600 800 254720
rect 0 253512 800 253632
rect 0 252288 800 252408
rect 0 251064 800 251184
rect 0 249840 800 249960
rect 0 248616 800 248736
rect 0 247392 800 247512
rect 0 246168 800 246288
rect 0 244944 800 245064
rect 0 243720 800 243840
rect 0 242496 800 242616
rect 0 241272 800 241392
rect 0 240048 800 240168
rect 0 238824 800 238944
rect 0 237600 800 237720
rect 0 236376 800 236496
rect 0 235152 800 235272
rect 0 233928 800 234048
rect 0 232840 800 232960
rect 0 231616 800 231736
rect 0 230392 800 230512
rect 0 229168 800 229288
rect 0 227944 800 228064
rect 0 226720 800 226840
rect 0 225496 800 225616
rect 0 224272 800 224392
rect 0 223048 800 223168
rect 0 221824 800 221944
rect 0 220600 800 220720
rect 0 219376 800 219496
rect 0 218152 800 218272
rect 0 216928 800 217048
rect 0 215704 800 215824
rect 0 214480 800 214600
rect 0 213256 800 213376
rect 0 212168 800 212288
rect 0 210944 800 211064
rect 0 209720 800 209840
rect 0 208496 800 208616
rect 0 207272 800 207392
rect 0 206048 800 206168
rect 0 204824 800 204944
rect 0 203600 800 203720
rect 0 202376 800 202496
rect 0 201152 800 201272
rect 0 199928 800 200048
rect 0 198704 800 198824
rect 0 197480 800 197600
rect 0 196256 800 196376
rect 0 195032 800 195152
rect 0 193808 800 193928
rect 0 192584 800 192704
rect 0 191360 800 191480
rect 0 190272 800 190392
rect 0 189048 800 189168
rect 0 187824 800 187944
rect 0 186600 800 186720
rect 0 185376 800 185496
rect 0 184152 800 184272
rect 0 182928 800 183048
rect 0 181704 800 181824
rect 0 180480 800 180600
rect 0 179256 800 179376
rect 0 178032 800 178152
rect 0 176808 800 176928
rect 0 175584 800 175704
rect 0 174360 800 174480
rect 0 173136 800 173256
rect 0 171912 800 172032
rect 0 170688 800 170808
rect 0 169600 800 169720
rect 0 168376 800 168496
rect 0 167152 800 167272
rect 0 165928 800 166048
rect 0 164704 800 164824
rect 0 163480 800 163600
rect 0 162256 800 162376
rect 0 161032 800 161152
rect 0 159808 800 159928
rect 0 158584 800 158704
rect 0 157360 800 157480
rect 0 156136 800 156256
rect 0 154912 800 155032
rect 0 153688 800 153808
rect 0 152464 800 152584
rect 0 151240 800 151360
rect 0 150016 800 150136
rect 0 148792 800 148912
rect 0 147704 800 147824
rect 0 146480 800 146600
rect 0 145256 800 145376
rect 0 144032 800 144152
rect 0 142808 800 142928
rect 0 141584 800 141704
rect 0 140360 800 140480
rect 0 139136 800 139256
rect 0 137912 800 138032
rect 0 136688 800 136808
rect 0 135464 800 135584
rect 0 134240 800 134360
rect 0 133016 800 133136
rect 0 131792 800 131912
rect 0 130568 800 130688
rect 0 129344 800 129464
rect 0 128120 800 128240
rect 0 127032 800 127152
rect 0 125808 800 125928
rect 0 124584 800 124704
rect 0 123360 800 123480
rect 0 122136 800 122256
rect 0 120912 800 121032
rect 0 119688 800 119808
rect 0 118464 800 118584
rect 0 117240 800 117360
rect 0 116016 800 116136
rect 0 114792 800 114912
rect 0 113568 800 113688
rect 0 112344 800 112464
rect 0 111120 800 111240
rect 0 109896 800 110016
rect 0 108672 800 108792
rect 0 107448 800 107568
rect 0 106360 800 106480
rect 0 105136 800 105256
rect 0 103912 800 104032
rect 0 102688 800 102808
rect 0 101464 800 101584
rect 0 100240 800 100360
rect 0 99016 800 99136
rect 0 97792 800 97912
rect 0 96568 800 96688
rect 0 95344 800 95464
rect 0 94120 800 94240
rect 0 92896 800 93016
rect 0 91672 800 91792
rect 0 90448 800 90568
rect 0 89224 800 89344
rect 0 88000 800 88120
rect 0 86776 800 86896
rect 0 85552 800 85672
rect 0 84464 800 84584
rect 0 83240 800 83360
rect 0 82016 800 82136
rect 0 80792 800 80912
rect 0 79568 800 79688
rect 0 78344 800 78464
rect 0 77120 800 77240
rect 0 75896 800 76016
rect 0 74672 800 74792
rect 0 73448 800 73568
rect 0 72224 800 72344
rect 0 71000 800 71120
rect 0 69776 800 69896
rect 0 68552 800 68672
rect 0 67328 800 67448
rect 0 66104 800 66224
rect 0 64880 800 65000
rect 0 63792 800 63912
rect 0 62568 800 62688
rect 0 61344 800 61464
rect 0 60120 800 60240
rect 0 58896 800 59016
rect 0 57672 800 57792
rect 0 56448 800 56568
rect 0 55224 800 55344
rect 0 54000 800 54120
rect 0 52776 800 52896
rect 0 51552 800 51672
rect 0 50328 800 50448
rect 0 49104 800 49224
rect 0 47880 800 48000
rect 0 46656 800 46776
rect 0 45432 800 45552
rect 0 44208 800 44328
rect 0 42984 800 43104
rect 0 41896 800 42016
rect 0 40672 800 40792
rect 0 39448 800 39568
rect 0 38224 800 38344
rect 0 37000 800 37120
rect 0 35776 800 35896
rect 0 34552 800 34672
rect 0 33328 800 33448
rect 0 32104 800 32224
rect 0 30880 800 31000
rect 0 29656 800 29776
rect 0 28432 800 28552
rect 0 27208 800 27328
rect 0 25984 800 26104
rect 0 24760 800 24880
rect 0 23536 800 23656
rect 0 22312 800 22432
rect 0 21224 800 21344
rect 0 20000 800 20120
rect 0 18776 800 18896
rect 0 17552 800 17672
rect 0 16328 800 16448
rect 0 15104 800 15224
rect 0 13880 800 14000
rect 0 12656 800 12776
rect 0 11432 800 11552
rect 0 10208 800 10328
rect 0 8984 800 9104
rect 0 7760 800 7880
rect 0 6536 800 6656
rect 0 5312 800 5432
rect 0 4088 800 4208
rect 0 2864 800 2984
rect 0 1640 800 1760
rect 0 552 800 672
<< obsm3 >>
rect 880 359240 234928 359413
rect 800 358296 234928 359240
rect 880 358016 234928 358296
rect 800 357072 234928 358016
rect 880 356792 234928 357072
rect 800 355848 234928 356792
rect 880 355568 234928 355848
rect 800 354624 234928 355568
rect 880 354344 234928 354624
rect 800 353400 234928 354344
rect 880 353120 234928 353400
rect 800 352176 234928 353120
rect 880 351896 234928 352176
rect 800 350952 234928 351896
rect 880 350672 234928 350952
rect 800 349728 234928 350672
rect 880 349448 234928 349728
rect 800 348504 234928 349448
rect 880 348224 234928 348504
rect 800 347280 234928 348224
rect 880 347000 234928 347280
rect 800 346056 234928 347000
rect 880 345776 234928 346056
rect 800 344832 234928 345776
rect 880 344552 234928 344832
rect 800 343608 234928 344552
rect 880 343328 234928 343608
rect 800 342384 234928 343328
rect 880 342104 234928 342384
rect 800 341160 234928 342104
rect 880 340880 234928 341160
rect 800 339936 234928 340880
rect 880 339656 234928 339936
rect 800 338848 234928 339656
rect 880 338568 234928 338848
rect 800 337624 234928 338568
rect 880 337344 234928 337624
rect 800 336400 234928 337344
rect 880 336120 234928 336400
rect 800 335176 234928 336120
rect 880 334896 234928 335176
rect 800 333952 234928 334896
rect 880 333672 234928 333952
rect 800 332728 234928 333672
rect 880 332448 234928 332728
rect 800 331504 234928 332448
rect 880 331224 234928 331504
rect 800 330280 234928 331224
rect 880 330000 234928 330280
rect 800 329056 234928 330000
rect 880 328776 234928 329056
rect 800 327832 234928 328776
rect 880 327552 234928 327832
rect 800 326608 234928 327552
rect 880 326328 234928 326608
rect 800 325384 234928 326328
rect 880 325104 234928 325384
rect 800 324160 234928 325104
rect 880 323880 234928 324160
rect 800 322936 234928 323880
rect 880 322656 234928 322936
rect 800 321712 234928 322656
rect 880 321432 234928 321712
rect 800 320488 234928 321432
rect 880 320208 234928 320488
rect 800 319264 234928 320208
rect 880 318984 234928 319264
rect 800 318176 234928 318984
rect 880 317896 234928 318176
rect 800 316952 234928 317896
rect 880 316672 234928 316952
rect 800 315728 234928 316672
rect 880 315448 234928 315728
rect 800 314504 234928 315448
rect 880 314224 234928 314504
rect 800 313280 234928 314224
rect 880 313000 234928 313280
rect 800 312056 234928 313000
rect 880 311776 234928 312056
rect 800 310832 234928 311776
rect 880 310552 234928 310832
rect 800 309608 234928 310552
rect 880 309328 234928 309608
rect 800 308384 234928 309328
rect 880 308104 234928 308384
rect 800 307160 234928 308104
rect 880 306880 234928 307160
rect 800 305936 234928 306880
rect 880 305656 234928 305936
rect 800 304712 234928 305656
rect 880 304432 234928 304712
rect 800 303488 234928 304432
rect 880 303208 234928 303488
rect 800 302264 234928 303208
rect 880 301984 234928 302264
rect 800 301040 234928 301984
rect 880 300760 234928 301040
rect 800 299816 234928 300760
rect 880 299536 234928 299816
rect 800 298592 234928 299536
rect 880 298312 234928 298592
rect 800 297368 234928 298312
rect 880 297088 234928 297368
rect 800 296280 234928 297088
rect 880 296000 234928 296280
rect 800 295056 234928 296000
rect 880 294776 234928 295056
rect 800 293832 234928 294776
rect 880 293552 234928 293832
rect 800 292608 234928 293552
rect 880 292328 234928 292608
rect 800 291384 234928 292328
rect 880 291104 234928 291384
rect 800 290160 234928 291104
rect 880 289880 234928 290160
rect 800 288936 234928 289880
rect 880 288656 234928 288936
rect 800 287712 234928 288656
rect 880 287432 234928 287712
rect 800 286488 234928 287432
rect 880 286208 234928 286488
rect 800 285264 234928 286208
rect 880 284984 234928 285264
rect 800 284040 234928 284984
rect 880 283760 234928 284040
rect 800 282816 234928 283760
rect 880 282536 234928 282816
rect 800 281592 234928 282536
rect 880 281312 234928 281592
rect 800 280368 234928 281312
rect 880 280088 234928 280368
rect 800 279144 234928 280088
rect 880 278864 234928 279144
rect 800 277920 234928 278864
rect 880 277640 234928 277920
rect 800 276696 234928 277640
rect 880 276416 234928 276696
rect 800 275608 234928 276416
rect 880 275328 234928 275608
rect 800 274384 234928 275328
rect 880 274104 234928 274384
rect 800 273160 234928 274104
rect 880 272880 234928 273160
rect 800 271936 234928 272880
rect 880 271656 234928 271936
rect 800 270712 234928 271656
rect 880 270432 234928 270712
rect 800 269488 234928 270432
rect 880 269208 234928 269488
rect 800 268264 234928 269208
rect 880 267984 234928 268264
rect 800 267040 234928 267984
rect 880 266760 234928 267040
rect 800 265816 234928 266760
rect 880 265536 234928 265816
rect 800 264592 234928 265536
rect 880 264312 234928 264592
rect 800 263368 234928 264312
rect 880 263088 234928 263368
rect 800 262144 234928 263088
rect 880 261864 234928 262144
rect 800 260920 234928 261864
rect 880 260640 234928 260920
rect 800 259696 234928 260640
rect 880 259416 234928 259696
rect 800 258472 234928 259416
rect 880 258192 234928 258472
rect 800 257248 234928 258192
rect 880 256968 234928 257248
rect 800 256024 234928 256968
rect 880 255744 234928 256024
rect 800 254800 234928 255744
rect 880 254520 234928 254800
rect 800 253712 234928 254520
rect 880 253432 234928 253712
rect 800 252488 234928 253432
rect 880 252208 234928 252488
rect 800 251264 234928 252208
rect 880 250984 234928 251264
rect 800 250040 234928 250984
rect 880 249760 234928 250040
rect 800 248816 234928 249760
rect 880 248536 234928 248816
rect 800 247592 234928 248536
rect 880 247312 234928 247592
rect 800 246368 234928 247312
rect 880 246088 234928 246368
rect 800 245144 234928 246088
rect 880 244864 234928 245144
rect 800 243920 234928 244864
rect 880 243640 234928 243920
rect 800 242696 234928 243640
rect 880 242416 234928 242696
rect 800 241472 234928 242416
rect 880 241192 234928 241472
rect 800 240248 234928 241192
rect 880 239968 234928 240248
rect 800 239024 234928 239968
rect 880 238744 234928 239024
rect 800 237800 234928 238744
rect 880 237520 234928 237800
rect 800 236576 234928 237520
rect 880 236296 234928 236576
rect 800 235352 234928 236296
rect 880 235072 234928 235352
rect 800 234128 234928 235072
rect 880 233848 234928 234128
rect 800 233040 234928 233848
rect 880 232760 234928 233040
rect 800 231816 234928 232760
rect 880 231536 234928 231816
rect 800 230592 234928 231536
rect 880 230312 234928 230592
rect 800 229368 234928 230312
rect 880 229088 234928 229368
rect 800 228144 234928 229088
rect 880 227864 234928 228144
rect 800 226920 234928 227864
rect 880 226640 234928 226920
rect 800 225696 234928 226640
rect 880 225416 234928 225696
rect 800 224472 234928 225416
rect 880 224192 234928 224472
rect 800 223248 234928 224192
rect 880 222968 234928 223248
rect 800 222024 234928 222968
rect 880 221744 234928 222024
rect 800 220800 234928 221744
rect 880 220520 234928 220800
rect 800 219576 234928 220520
rect 880 219296 234928 219576
rect 800 218352 234928 219296
rect 880 218072 234928 218352
rect 800 217128 234928 218072
rect 880 216848 234928 217128
rect 800 215904 234928 216848
rect 880 215624 234928 215904
rect 800 214680 234928 215624
rect 880 214400 234928 214680
rect 800 213456 234928 214400
rect 880 213176 234928 213456
rect 800 212368 234928 213176
rect 880 212088 234928 212368
rect 800 211144 234928 212088
rect 880 210864 234928 211144
rect 800 209920 234928 210864
rect 880 209640 234928 209920
rect 800 208696 234928 209640
rect 880 208416 234928 208696
rect 800 207472 234928 208416
rect 880 207192 234928 207472
rect 800 206248 234928 207192
rect 880 205968 234928 206248
rect 800 205024 234928 205968
rect 880 204744 234928 205024
rect 800 203800 234928 204744
rect 880 203520 234928 203800
rect 800 202576 234928 203520
rect 880 202296 234928 202576
rect 800 201352 234928 202296
rect 880 201072 234928 201352
rect 800 200128 234928 201072
rect 880 199848 234928 200128
rect 800 198904 234928 199848
rect 880 198624 234928 198904
rect 800 197680 234928 198624
rect 880 197400 234928 197680
rect 800 196456 234928 197400
rect 880 196176 234928 196456
rect 800 195232 234928 196176
rect 880 194952 234928 195232
rect 800 194008 234928 194952
rect 880 193728 234928 194008
rect 800 192784 234928 193728
rect 880 192504 234928 192784
rect 800 191560 234928 192504
rect 880 191280 234928 191560
rect 800 190472 234928 191280
rect 880 190192 234928 190472
rect 800 189248 234928 190192
rect 880 188968 234928 189248
rect 800 188024 234928 188968
rect 880 187744 234928 188024
rect 800 186800 234928 187744
rect 880 186520 234928 186800
rect 800 185576 234928 186520
rect 880 185296 234928 185576
rect 800 184352 234928 185296
rect 880 184072 234928 184352
rect 800 183128 234928 184072
rect 880 182848 234928 183128
rect 800 181904 234928 182848
rect 880 181624 234928 181904
rect 800 180680 234928 181624
rect 880 180400 234928 180680
rect 800 179456 234928 180400
rect 880 179176 234928 179456
rect 800 178232 234928 179176
rect 880 177952 234928 178232
rect 800 177008 234928 177952
rect 880 176728 234928 177008
rect 800 175784 234928 176728
rect 880 175504 234928 175784
rect 800 174560 234928 175504
rect 880 174280 234928 174560
rect 800 173336 234928 174280
rect 880 173056 234928 173336
rect 800 172112 234928 173056
rect 880 171832 234928 172112
rect 800 170888 234928 171832
rect 880 170608 234928 170888
rect 800 169800 234928 170608
rect 880 169520 234928 169800
rect 800 168576 234928 169520
rect 880 168296 234928 168576
rect 800 167352 234928 168296
rect 880 167072 234928 167352
rect 800 166128 234928 167072
rect 880 165848 234928 166128
rect 800 164904 234928 165848
rect 880 164624 234928 164904
rect 800 163680 234928 164624
rect 880 163400 234928 163680
rect 800 162456 234928 163400
rect 880 162176 234928 162456
rect 800 161232 234928 162176
rect 880 160952 234928 161232
rect 800 160008 234928 160952
rect 880 159728 234928 160008
rect 800 158784 234928 159728
rect 880 158504 234928 158784
rect 800 157560 234928 158504
rect 880 157280 234928 157560
rect 800 156336 234928 157280
rect 880 156056 234928 156336
rect 800 155112 234928 156056
rect 880 154832 234928 155112
rect 800 153888 234928 154832
rect 880 153608 234928 153888
rect 800 152664 234928 153608
rect 880 152384 234928 152664
rect 800 151440 234928 152384
rect 880 151160 234928 151440
rect 800 150216 234928 151160
rect 880 149936 234928 150216
rect 800 148992 234928 149936
rect 880 148712 234928 148992
rect 800 147904 234928 148712
rect 880 147624 234928 147904
rect 800 146680 234928 147624
rect 880 146400 234928 146680
rect 800 145456 234928 146400
rect 880 145176 234928 145456
rect 800 144232 234928 145176
rect 880 143952 234928 144232
rect 800 143008 234928 143952
rect 880 142728 234928 143008
rect 800 141784 234928 142728
rect 880 141504 234928 141784
rect 800 140560 234928 141504
rect 880 140280 234928 140560
rect 800 139336 234928 140280
rect 880 139056 234928 139336
rect 800 138112 234928 139056
rect 880 137832 234928 138112
rect 800 136888 234928 137832
rect 880 136608 234928 136888
rect 800 135664 234928 136608
rect 880 135384 234928 135664
rect 800 134440 234928 135384
rect 880 134160 234928 134440
rect 800 133216 234928 134160
rect 880 132936 234928 133216
rect 800 131992 234928 132936
rect 880 131712 234928 131992
rect 800 130768 234928 131712
rect 880 130488 234928 130768
rect 800 129544 234928 130488
rect 880 129264 234928 129544
rect 800 128320 234928 129264
rect 880 128040 234928 128320
rect 800 127232 234928 128040
rect 880 126952 234928 127232
rect 800 126008 234928 126952
rect 880 125728 234928 126008
rect 800 124784 234928 125728
rect 880 124504 234928 124784
rect 800 123560 234928 124504
rect 880 123280 234928 123560
rect 800 122336 234928 123280
rect 880 122056 234928 122336
rect 800 121112 234928 122056
rect 880 120832 234928 121112
rect 800 119888 234928 120832
rect 880 119608 234928 119888
rect 800 118664 234928 119608
rect 880 118384 234928 118664
rect 800 117440 234928 118384
rect 880 117160 234928 117440
rect 800 116216 234928 117160
rect 880 115936 234928 116216
rect 800 114992 234928 115936
rect 880 114712 234928 114992
rect 800 113768 234928 114712
rect 880 113488 234928 113768
rect 800 112544 234928 113488
rect 880 112264 234928 112544
rect 800 111320 234928 112264
rect 880 111040 234928 111320
rect 800 110096 234928 111040
rect 880 109816 234928 110096
rect 800 108872 234928 109816
rect 880 108592 234928 108872
rect 800 107648 234928 108592
rect 880 107368 234928 107648
rect 800 106560 234928 107368
rect 880 106280 234928 106560
rect 800 105336 234928 106280
rect 880 105056 234928 105336
rect 800 104112 234928 105056
rect 880 103832 234928 104112
rect 800 102888 234928 103832
rect 880 102608 234928 102888
rect 800 101664 234928 102608
rect 880 101384 234928 101664
rect 800 100440 234928 101384
rect 880 100160 234928 100440
rect 800 99216 234928 100160
rect 880 98936 234928 99216
rect 800 97992 234928 98936
rect 880 97712 234928 97992
rect 800 96768 234928 97712
rect 880 96488 234928 96768
rect 800 95544 234928 96488
rect 880 95264 234928 95544
rect 800 94320 234928 95264
rect 880 94040 234928 94320
rect 800 93096 234928 94040
rect 880 92816 234928 93096
rect 800 91872 234928 92816
rect 880 91592 234928 91872
rect 800 90648 234928 91592
rect 880 90368 234928 90648
rect 800 89424 234928 90368
rect 880 89144 234928 89424
rect 800 88200 234928 89144
rect 880 87920 234928 88200
rect 800 86976 234928 87920
rect 880 86696 234928 86976
rect 800 85752 234928 86696
rect 880 85472 234928 85752
rect 800 84664 234928 85472
rect 880 84384 234928 84664
rect 800 83440 234928 84384
rect 880 83160 234928 83440
rect 800 82216 234928 83160
rect 880 81936 234928 82216
rect 800 80992 234928 81936
rect 880 80712 234928 80992
rect 800 79768 234928 80712
rect 880 79488 234928 79768
rect 800 78544 234928 79488
rect 880 78264 234928 78544
rect 800 77320 234928 78264
rect 880 77040 234928 77320
rect 800 76096 234928 77040
rect 880 75816 234928 76096
rect 800 74872 234928 75816
rect 880 74592 234928 74872
rect 800 73648 234928 74592
rect 880 73368 234928 73648
rect 800 72424 234928 73368
rect 880 72144 234928 72424
rect 800 71200 234928 72144
rect 880 70920 234928 71200
rect 800 69976 234928 70920
rect 880 69696 234928 69976
rect 800 68752 234928 69696
rect 880 68472 234928 68752
rect 800 67528 234928 68472
rect 880 67248 234928 67528
rect 800 66304 234928 67248
rect 880 66024 234928 66304
rect 800 65080 234928 66024
rect 880 64800 234928 65080
rect 800 63992 234928 64800
rect 880 63712 234928 63992
rect 800 62768 234928 63712
rect 880 62488 234928 62768
rect 800 61544 234928 62488
rect 880 61264 234928 61544
rect 800 60320 234928 61264
rect 880 60040 234928 60320
rect 800 59096 234928 60040
rect 880 58816 234928 59096
rect 800 57872 234928 58816
rect 880 57592 234928 57872
rect 800 56648 234928 57592
rect 880 56368 234928 56648
rect 800 55424 234928 56368
rect 880 55144 234928 55424
rect 800 54200 234928 55144
rect 880 53920 234928 54200
rect 800 52976 234928 53920
rect 880 52696 234928 52976
rect 800 51752 234928 52696
rect 880 51472 234928 51752
rect 800 50528 234928 51472
rect 880 50248 234928 50528
rect 800 49304 234928 50248
rect 880 49024 234928 49304
rect 800 48080 234928 49024
rect 880 47800 234928 48080
rect 800 46856 234928 47800
rect 880 46576 234928 46856
rect 800 45632 234928 46576
rect 880 45352 234928 45632
rect 800 44408 234928 45352
rect 880 44128 234928 44408
rect 800 43184 234928 44128
rect 880 42904 234928 43184
rect 800 42096 234928 42904
rect 880 41816 234928 42096
rect 800 40872 234928 41816
rect 880 40592 234928 40872
rect 800 39648 234928 40592
rect 880 39368 234928 39648
rect 800 38424 234928 39368
rect 880 38144 234928 38424
rect 800 37200 234928 38144
rect 880 36920 234928 37200
rect 800 35976 234928 36920
rect 880 35696 234928 35976
rect 800 34752 234928 35696
rect 880 34472 234928 34752
rect 800 33528 234928 34472
rect 880 33248 234928 33528
rect 800 32304 234928 33248
rect 880 32024 234928 32304
rect 800 31080 234928 32024
rect 880 30800 234928 31080
rect 800 29856 234928 30800
rect 880 29576 234928 29856
rect 800 28632 234928 29576
rect 880 28352 234928 28632
rect 800 27408 234928 28352
rect 880 27128 234928 27408
rect 800 26184 234928 27128
rect 880 25904 234928 26184
rect 800 24960 234928 25904
rect 880 24680 234928 24960
rect 800 23736 234928 24680
rect 880 23456 234928 23736
rect 800 22512 234928 23456
rect 880 22232 234928 22512
rect 800 21424 234928 22232
rect 880 21144 234928 21424
rect 800 20200 234928 21144
rect 880 19920 234928 20200
rect 800 18976 234928 19920
rect 880 18696 234928 18976
rect 800 17752 234928 18696
rect 880 17472 234928 17752
rect 800 16528 234928 17472
rect 880 16248 234928 16528
rect 800 15304 234928 16248
rect 880 15024 234928 15304
rect 800 14080 234928 15024
rect 880 13800 234928 14080
rect 800 12856 234928 13800
rect 880 12576 234928 12856
rect 800 11632 234928 12576
rect 880 11352 234928 11632
rect 800 10408 234928 11352
rect 880 10128 234928 10408
rect 800 9184 234928 10128
rect 880 8904 234928 9184
rect 800 7960 234928 8904
rect 880 7680 234928 7960
rect 800 6736 234928 7680
rect 880 6456 234928 6736
rect 800 5512 234928 6456
rect 880 5232 234928 5512
rect 800 4288 234928 5232
rect 880 4008 234928 4288
rect 800 3064 234928 4008
rect 880 2784 234928 3064
rect 800 1840 234928 2784
rect 880 1560 234928 1840
rect 800 752 234928 1560
rect 880 579 234928 752
<< metal4 >>
rect 4208 2128 4528 357456
rect 19568 2128 19888 357456
rect 34928 2128 35248 357456
rect 50288 2128 50608 357456
rect 65648 2128 65968 357456
rect 81008 2128 81328 357456
rect 96368 2128 96688 357456
rect 111728 2128 112048 357456
rect 127088 2128 127408 357456
rect 142448 2128 142768 357456
rect 157808 2128 158128 357456
rect 173168 2128 173488 357456
rect 188528 2128 188848 357456
rect 203888 2128 204208 357456
rect 219248 2128 219568 357456
rect 234608 2128 234928 357456
<< obsm4 >>
rect 1531 2347 4128 350981
rect 4608 2347 19488 350981
rect 19968 2347 34848 350981
rect 35328 2347 50208 350981
rect 50688 2347 65568 350981
rect 66048 2347 80928 350981
rect 81408 2347 96288 350981
rect 96768 2347 111648 350981
rect 112128 2347 127008 350981
rect 127488 2347 142368 350981
rect 142848 2347 157728 350981
rect 158208 2347 163517 350981
<< labels >>
rlabel metal3 s 0 161032 800 161152 6 bb_addr0[0]
port 1 nsew signal output
rlabel metal3 s 0 226720 800 226840 6 bb_addr0[10]
port 2 nsew signal output
rlabel metal3 s 0 232840 800 232960 6 bb_addr0[11]
port 3 nsew signal output
rlabel metal3 s 0 238824 800 238944 6 bb_addr0[12]
port 4 nsew signal output
rlabel metal3 s 0 244944 800 245064 6 bb_addr0[13]
port 5 nsew signal output
rlabel metal3 s 0 251064 800 251184 6 bb_addr0[14]
port 6 nsew signal output
rlabel metal3 s 0 257048 800 257168 6 bb_addr0[15]
port 7 nsew signal output
rlabel metal3 s 0 263168 800 263288 6 bb_addr0[16]
port 8 nsew signal output
rlabel metal3 s 0 269288 800 269408 6 bb_addr0[17]
port 9 nsew signal output
rlabel metal3 s 0 275408 800 275528 6 bb_addr0[18]
port 10 nsew signal output
rlabel metal3 s 0 281392 800 281512 6 bb_addr0[19]
port 11 nsew signal output
rlabel metal3 s 0 168376 800 168496 6 bb_addr0[1]
port 12 nsew signal output
rlabel metal3 s 0 287512 800 287632 6 bb_addr0[20]
port 13 nsew signal output
rlabel metal3 s 0 293632 800 293752 6 bb_addr0[21]
port 14 nsew signal output
rlabel metal3 s 0 299616 800 299736 6 bb_addr0[22]
port 15 nsew signal output
rlabel metal3 s 0 305736 800 305856 6 bb_addr0[23]
port 16 nsew signal output
rlabel metal3 s 0 311856 800 311976 6 bb_addr0[24]
port 17 nsew signal output
rlabel metal3 s 0 317976 800 318096 6 bb_addr0[25]
port 18 nsew signal output
rlabel metal3 s 0 323960 800 324080 6 bb_addr0[26]
port 19 nsew signal output
rlabel metal3 s 0 330080 800 330200 6 bb_addr0[27]
port 20 nsew signal output
rlabel metal3 s 0 336200 800 336320 6 bb_addr0[28]
port 21 nsew signal output
rlabel metal3 s 0 342184 800 342304 6 bb_addr0[29]
port 22 nsew signal output
rlabel metal3 s 0 175584 800 175704 6 bb_addr0[2]
port 23 nsew signal output
rlabel metal3 s 0 348304 800 348424 6 bb_addr0[30]
port 24 nsew signal output
rlabel metal3 s 0 354424 800 354544 6 bb_addr0[31]
port 25 nsew signal output
rlabel metal3 s 0 182928 800 183048 6 bb_addr0[3]
port 26 nsew signal output
rlabel metal3 s 0 190272 800 190392 6 bb_addr0[4]
port 27 nsew signal output
rlabel metal3 s 0 196256 800 196376 6 bb_addr0[5]
port 28 nsew signal output
rlabel metal3 s 0 202376 800 202496 6 bb_addr0[6]
port 29 nsew signal output
rlabel metal3 s 0 208496 800 208616 6 bb_addr0[7]
port 30 nsew signal output
rlabel metal3 s 0 214480 800 214600 6 bb_addr0[8]
port 31 nsew signal output
rlabel metal3 s 0 220600 800 220720 6 bb_addr0[9]
port 32 nsew signal output
rlabel metal3 s 0 162256 800 162376 6 bb_addr1[0]
port 33 nsew signal output
rlabel metal3 s 0 227944 800 228064 6 bb_addr1[10]
port 34 nsew signal output
rlabel metal3 s 0 233928 800 234048 6 bb_addr1[11]
port 35 nsew signal output
rlabel metal3 s 0 240048 800 240168 6 bb_addr1[12]
port 36 nsew signal output
rlabel metal3 s 0 246168 800 246288 6 bb_addr1[13]
port 37 nsew signal output
rlabel metal3 s 0 252288 800 252408 6 bb_addr1[14]
port 38 nsew signal output
rlabel metal3 s 0 258272 800 258392 6 bb_addr1[15]
port 39 nsew signal output
rlabel metal3 s 0 264392 800 264512 6 bb_addr1[16]
port 40 nsew signal output
rlabel metal3 s 0 270512 800 270632 6 bb_addr1[17]
port 41 nsew signal output
rlabel metal3 s 0 276496 800 276616 6 bb_addr1[18]
port 42 nsew signal output
rlabel metal3 s 0 282616 800 282736 6 bb_addr1[19]
port 43 nsew signal output
rlabel metal3 s 0 169600 800 169720 6 bb_addr1[1]
port 44 nsew signal output
rlabel metal3 s 0 288736 800 288856 6 bb_addr1[20]
port 45 nsew signal output
rlabel metal3 s 0 294856 800 294976 6 bb_addr1[21]
port 46 nsew signal output
rlabel metal3 s 0 300840 800 300960 6 bb_addr1[22]
port 47 nsew signal output
rlabel metal3 s 0 306960 800 307080 6 bb_addr1[23]
port 48 nsew signal output
rlabel metal3 s 0 313080 800 313200 6 bb_addr1[24]
port 49 nsew signal output
rlabel metal3 s 0 319064 800 319184 6 bb_addr1[25]
port 50 nsew signal output
rlabel metal3 s 0 325184 800 325304 6 bb_addr1[26]
port 51 nsew signal output
rlabel metal3 s 0 331304 800 331424 6 bb_addr1[27]
port 52 nsew signal output
rlabel metal3 s 0 337424 800 337544 6 bb_addr1[28]
port 53 nsew signal output
rlabel metal3 s 0 343408 800 343528 6 bb_addr1[29]
port 54 nsew signal output
rlabel metal3 s 0 176808 800 176928 6 bb_addr1[2]
port 55 nsew signal output
rlabel metal3 s 0 349528 800 349648 6 bb_addr1[30]
port 56 nsew signal output
rlabel metal3 s 0 355648 800 355768 6 bb_addr1[31]
port 57 nsew signal output
rlabel metal3 s 0 184152 800 184272 6 bb_addr1[3]
port 58 nsew signal output
rlabel metal3 s 0 191360 800 191480 6 bb_addr1[4]
port 59 nsew signal output
rlabel metal3 s 0 197480 800 197600 6 bb_addr1[5]
port 60 nsew signal output
rlabel metal3 s 0 203600 800 203720 6 bb_addr1[6]
port 61 nsew signal output
rlabel metal3 s 0 209720 800 209840 6 bb_addr1[7]
port 62 nsew signal output
rlabel metal3 s 0 215704 800 215824 6 bb_addr1[8]
port 63 nsew signal output
rlabel metal3 s 0 221824 800 221944 6 bb_addr1[9]
port 64 nsew signal output
rlabel metal3 s 0 157360 800 157480 6 bb_csb0
port 65 nsew signal output
rlabel metal3 s 0 158584 800 158704 6 bb_csb1
port 66 nsew signal output
rlabel metal3 s 0 163480 800 163600 6 bb_din0[0]
port 67 nsew signal output
rlabel metal3 s 0 229168 800 229288 6 bb_din0[10]
port 68 nsew signal output
rlabel metal3 s 0 235152 800 235272 6 bb_din0[11]
port 69 nsew signal output
rlabel metal3 s 0 241272 800 241392 6 bb_din0[12]
port 70 nsew signal output
rlabel metal3 s 0 247392 800 247512 6 bb_din0[13]
port 71 nsew signal output
rlabel metal3 s 0 253512 800 253632 6 bb_din0[14]
port 72 nsew signal output
rlabel metal3 s 0 259496 800 259616 6 bb_din0[15]
port 73 nsew signal output
rlabel metal3 s 0 265616 800 265736 6 bb_din0[16]
port 74 nsew signal output
rlabel metal3 s 0 271736 800 271856 6 bb_din0[17]
port 75 nsew signal output
rlabel metal3 s 0 277720 800 277840 6 bb_din0[18]
port 76 nsew signal output
rlabel metal3 s 0 283840 800 283960 6 bb_din0[19]
port 77 nsew signal output
rlabel metal3 s 0 170688 800 170808 6 bb_din0[1]
port 78 nsew signal output
rlabel metal3 s 0 289960 800 290080 6 bb_din0[20]
port 79 nsew signal output
rlabel metal3 s 0 296080 800 296200 6 bb_din0[21]
port 80 nsew signal output
rlabel metal3 s 0 302064 800 302184 6 bb_din0[22]
port 81 nsew signal output
rlabel metal3 s 0 308184 800 308304 6 bb_din0[23]
port 82 nsew signal output
rlabel metal3 s 0 314304 800 314424 6 bb_din0[24]
port 83 nsew signal output
rlabel metal3 s 0 320288 800 320408 6 bb_din0[25]
port 84 nsew signal output
rlabel metal3 s 0 326408 800 326528 6 bb_din0[26]
port 85 nsew signal output
rlabel metal3 s 0 332528 800 332648 6 bb_din0[27]
port 86 nsew signal output
rlabel metal3 s 0 338648 800 338768 6 bb_din0[28]
port 87 nsew signal output
rlabel metal3 s 0 344632 800 344752 6 bb_din0[29]
port 88 nsew signal output
rlabel metal3 s 0 178032 800 178152 6 bb_din0[2]
port 89 nsew signal output
rlabel metal3 s 0 350752 800 350872 6 bb_din0[30]
port 90 nsew signal output
rlabel metal3 s 0 356872 800 356992 6 bb_din0[31]
port 91 nsew signal output
rlabel metal3 s 0 185376 800 185496 6 bb_din0[3]
port 92 nsew signal output
rlabel metal3 s 0 192584 800 192704 6 bb_din0[4]
port 93 nsew signal output
rlabel metal3 s 0 198704 800 198824 6 bb_din0[5]
port 94 nsew signal output
rlabel metal3 s 0 204824 800 204944 6 bb_din0[6]
port 95 nsew signal output
rlabel metal3 s 0 210944 800 211064 6 bb_din0[7]
port 96 nsew signal output
rlabel metal3 s 0 216928 800 217048 6 bb_din0[8]
port 97 nsew signal output
rlabel metal3 s 0 223048 800 223168 6 bb_din0[9]
port 98 nsew signal output
rlabel metal3 s 0 164704 800 164824 6 bb_dout0[0]
port 99 nsew signal input
rlabel metal3 s 0 230392 800 230512 6 bb_dout0[10]
port 100 nsew signal input
rlabel metal3 s 0 236376 800 236496 6 bb_dout0[11]
port 101 nsew signal input
rlabel metal3 s 0 242496 800 242616 6 bb_dout0[12]
port 102 nsew signal input
rlabel metal3 s 0 248616 800 248736 6 bb_dout0[13]
port 103 nsew signal input
rlabel metal3 s 0 254600 800 254720 6 bb_dout0[14]
port 104 nsew signal input
rlabel metal3 s 0 260720 800 260840 6 bb_dout0[15]
port 105 nsew signal input
rlabel metal3 s 0 266840 800 266960 6 bb_dout0[16]
port 106 nsew signal input
rlabel metal3 s 0 272960 800 273080 6 bb_dout0[17]
port 107 nsew signal input
rlabel metal3 s 0 278944 800 279064 6 bb_dout0[18]
port 108 nsew signal input
rlabel metal3 s 0 285064 800 285184 6 bb_dout0[19]
port 109 nsew signal input
rlabel metal3 s 0 171912 800 172032 6 bb_dout0[1]
port 110 nsew signal input
rlabel metal3 s 0 291184 800 291304 6 bb_dout0[20]
port 111 nsew signal input
rlabel metal3 s 0 297168 800 297288 6 bb_dout0[21]
port 112 nsew signal input
rlabel metal3 s 0 303288 800 303408 6 bb_dout0[22]
port 113 nsew signal input
rlabel metal3 s 0 309408 800 309528 6 bb_dout0[23]
port 114 nsew signal input
rlabel metal3 s 0 315528 800 315648 6 bb_dout0[24]
port 115 nsew signal input
rlabel metal3 s 0 321512 800 321632 6 bb_dout0[25]
port 116 nsew signal input
rlabel metal3 s 0 327632 800 327752 6 bb_dout0[26]
port 117 nsew signal input
rlabel metal3 s 0 333752 800 333872 6 bb_dout0[27]
port 118 nsew signal input
rlabel metal3 s 0 339736 800 339856 6 bb_dout0[28]
port 119 nsew signal input
rlabel metal3 s 0 345856 800 345976 6 bb_dout0[29]
port 120 nsew signal input
rlabel metal3 s 0 179256 800 179376 6 bb_dout0[2]
port 121 nsew signal input
rlabel metal3 s 0 351976 800 352096 6 bb_dout0[30]
port 122 nsew signal input
rlabel metal3 s 0 358096 800 358216 6 bb_dout0[31]
port 123 nsew signal input
rlabel metal3 s 0 186600 800 186720 6 bb_dout0[3]
port 124 nsew signal input
rlabel metal3 s 0 193808 800 193928 6 bb_dout0[4]
port 125 nsew signal input
rlabel metal3 s 0 199928 800 200048 6 bb_dout0[5]
port 126 nsew signal input
rlabel metal3 s 0 206048 800 206168 6 bb_dout0[6]
port 127 nsew signal input
rlabel metal3 s 0 212168 800 212288 6 bb_dout0[7]
port 128 nsew signal input
rlabel metal3 s 0 218152 800 218272 6 bb_dout0[8]
port 129 nsew signal input
rlabel metal3 s 0 224272 800 224392 6 bb_dout0[9]
port 130 nsew signal input
rlabel metal3 s 0 165928 800 166048 6 bb_dout1[0]
port 131 nsew signal input
rlabel metal3 s 0 231616 800 231736 6 bb_dout1[10]
port 132 nsew signal input
rlabel metal3 s 0 237600 800 237720 6 bb_dout1[11]
port 133 nsew signal input
rlabel metal3 s 0 243720 800 243840 6 bb_dout1[12]
port 134 nsew signal input
rlabel metal3 s 0 249840 800 249960 6 bb_dout1[13]
port 135 nsew signal input
rlabel metal3 s 0 255824 800 255944 6 bb_dout1[14]
port 136 nsew signal input
rlabel metal3 s 0 261944 800 262064 6 bb_dout1[15]
port 137 nsew signal input
rlabel metal3 s 0 268064 800 268184 6 bb_dout1[16]
port 138 nsew signal input
rlabel metal3 s 0 274184 800 274304 6 bb_dout1[17]
port 139 nsew signal input
rlabel metal3 s 0 280168 800 280288 6 bb_dout1[18]
port 140 nsew signal input
rlabel metal3 s 0 286288 800 286408 6 bb_dout1[19]
port 141 nsew signal input
rlabel metal3 s 0 173136 800 173256 6 bb_dout1[1]
port 142 nsew signal input
rlabel metal3 s 0 292408 800 292528 6 bb_dout1[20]
port 143 nsew signal input
rlabel metal3 s 0 298392 800 298512 6 bb_dout1[21]
port 144 nsew signal input
rlabel metal3 s 0 304512 800 304632 6 bb_dout1[22]
port 145 nsew signal input
rlabel metal3 s 0 310632 800 310752 6 bb_dout1[23]
port 146 nsew signal input
rlabel metal3 s 0 316752 800 316872 6 bb_dout1[24]
port 147 nsew signal input
rlabel metal3 s 0 322736 800 322856 6 bb_dout1[25]
port 148 nsew signal input
rlabel metal3 s 0 328856 800 328976 6 bb_dout1[26]
port 149 nsew signal input
rlabel metal3 s 0 334976 800 335096 6 bb_dout1[27]
port 150 nsew signal input
rlabel metal3 s 0 340960 800 341080 6 bb_dout1[28]
port 151 nsew signal input
rlabel metal3 s 0 347080 800 347200 6 bb_dout1[29]
port 152 nsew signal input
rlabel metal3 s 0 180480 800 180600 6 bb_dout1[2]
port 153 nsew signal input
rlabel metal3 s 0 353200 800 353320 6 bb_dout1[30]
port 154 nsew signal input
rlabel metal3 s 0 359320 800 359440 6 bb_dout1[31]
port 155 nsew signal input
rlabel metal3 s 0 187824 800 187944 6 bb_dout1[3]
port 156 nsew signal input
rlabel metal3 s 0 195032 800 195152 6 bb_dout1[4]
port 157 nsew signal input
rlabel metal3 s 0 201152 800 201272 6 bb_dout1[5]
port 158 nsew signal input
rlabel metal3 s 0 207272 800 207392 6 bb_dout1[6]
port 159 nsew signal input
rlabel metal3 s 0 213256 800 213376 6 bb_dout1[7]
port 160 nsew signal input
rlabel metal3 s 0 219376 800 219496 6 bb_dout1[8]
port 161 nsew signal input
rlabel metal3 s 0 225496 800 225616 6 bb_dout1[9]
port 162 nsew signal input
rlabel metal3 s 0 159808 800 159928 6 bb_web0
port 163 nsew signal output
rlabel metal3 s 0 167152 800 167272 6 bb_wmask0[0]
port 164 nsew signal output
rlabel metal3 s 0 174360 800 174480 6 bb_wmask0[1]
port 165 nsew signal output
rlabel metal3 s 0 181704 800 181824 6 bb_wmask0[2]
port 166 nsew signal output
rlabel metal3 s 0 189048 800 189168 6 bb_wmask0[3]
port 167 nsew signal output
rlabel metal2 s 1582 0 1638 800 6 clk_g
port 168 nsew signal input
rlabel metal2 s 14370 0 14426 800 6 io_gecerli
port 169 nsew signal output
rlabel metal2 s 17498 0 17554 800 6 io_oeb[0]
port 170 nsew signal output
rlabel metal2 s 81530 0 81586 800 6 io_oeb[10]
port 171 nsew signal output
rlabel metal2 s 87970 0 88026 800 6 io_oeb[11]
port 172 nsew signal output
rlabel metal2 s 94318 0 94374 800 6 io_oeb[12]
port 173 nsew signal output
rlabel metal2 s 100758 0 100814 800 6 io_oeb[13]
port 174 nsew signal output
rlabel metal2 s 107106 0 107162 800 6 io_oeb[14]
port 175 nsew signal output
rlabel metal2 s 113546 0 113602 800 6 io_oeb[15]
port 176 nsew signal output
rlabel metal2 s 119986 0 120042 800 6 io_oeb[16]
port 177 nsew signal output
rlabel metal2 s 126334 0 126390 800 6 io_oeb[17]
port 178 nsew signal output
rlabel metal2 s 132774 0 132830 800 6 io_oeb[18]
port 179 nsew signal output
rlabel metal2 s 139122 0 139178 800 6 io_oeb[19]
port 180 nsew signal output
rlabel metal2 s 23938 0 23994 800 6 io_oeb[1]
port 181 nsew signal output
rlabel metal2 s 145562 0 145618 800 6 io_oeb[20]
port 182 nsew signal output
rlabel metal2 s 151910 0 151966 800 6 io_oeb[21]
port 183 nsew signal output
rlabel metal2 s 158350 0 158406 800 6 io_oeb[22]
port 184 nsew signal output
rlabel metal2 s 164790 0 164846 800 6 io_oeb[23]
port 185 nsew signal output
rlabel metal2 s 171138 0 171194 800 6 io_oeb[24]
port 186 nsew signal output
rlabel metal2 s 177578 0 177634 800 6 io_oeb[25]
port 187 nsew signal output
rlabel metal2 s 183926 0 183982 800 6 io_oeb[26]
port 188 nsew signal output
rlabel metal2 s 190366 0 190422 800 6 io_oeb[27]
port 189 nsew signal output
rlabel metal2 s 196714 0 196770 800 6 io_oeb[28]
port 190 nsew signal output
rlabel metal2 s 203154 0 203210 800 6 io_oeb[29]
port 191 nsew signal output
rlabel metal2 s 30378 0 30434 800 6 io_oeb[2]
port 192 nsew signal output
rlabel metal2 s 209594 0 209650 800 6 io_oeb[30]
port 193 nsew signal output
rlabel metal2 s 215942 0 215998 800 6 io_oeb[31]
port 194 nsew signal output
rlabel metal2 s 222382 0 222438 800 6 io_oeb[32]
port 195 nsew signal output
rlabel metal2 s 225602 0 225658 800 6 io_oeb[33]
port 196 nsew signal output
rlabel metal2 s 228730 0 228786 800 6 io_oeb[34]
port 197 nsew signal output
rlabel metal2 s 231950 0 232006 800 6 io_oeb[35]
port 198 nsew signal output
rlabel metal2 s 235170 0 235226 800 6 io_oeb[36]
port 199 nsew signal output
rlabel metal2 s 238390 0 238446 800 6 io_oeb[37]
port 200 nsew signal output
rlabel metal2 s 36726 0 36782 800 6 io_oeb[3]
port 201 nsew signal output
rlabel metal2 s 43166 0 43222 800 6 io_oeb[4]
port 202 nsew signal output
rlabel metal2 s 49514 0 49570 800 6 io_oeb[5]
port 203 nsew signal output
rlabel metal2 s 55954 0 56010 800 6 io_oeb[6]
port 204 nsew signal output
rlabel metal2 s 62302 0 62358 800 6 io_oeb[7]
port 205 nsew signal output
rlabel metal2 s 68742 0 68798 800 6 io_oeb[8]
port 206 nsew signal output
rlabel metal2 s 75182 0 75238 800 6 io_oeb[9]
port 207 nsew signal output
rlabel metal2 s 20718 0 20774 800 6 io_ps[0]
port 208 nsew signal output
rlabel metal2 s 84750 0 84806 800 6 io_ps[10]
port 209 nsew signal output
rlabel metal2 s 91190 0 91246 800 6 io_ps[11]
port 210 nsew signal output
rlabel metal2 s 97538 0 97594 800 6 io_ps[12]
port 211 nsew signal output
rlabel metal2 s 103978 0 104034 800 6 io_ps[13]
port 212 nsew signal output
rlabel metal2 s 110326 0 110382 800 6 io_ps[14]
port 213 nsew signal output
rlabel metal2 s 116766 0 116822 800 6 io_ps[15]
port 214 nsew signal output
rlabel metal2 s 123114 0 123170 800 6 io_ps[16]
port 215 nsew signal output
rlabel metal2 s 129554 0 129610 800 6 io_ps[17]
port 216 nsew signal output
rlabel metal2 s 135994 0 136050 800 6 io_ps[18]
port 217 nsew signal output
rlabel metal2 s 142342 0 142398 800 6 io_ps[19]
port 218 nsew signal output
rlabel metal2 s 27158 0 27214 800 6 io_ps[1]
port 219 nsew signal output
rlabel metal2 s 148782 0 148838 800 6 io_ps[20]
port 220 nsew signal output
rlabel metal2 s 155130 0 155186 800 6 io_ps[21]
port 221 nsew signal output
rlabel metal2 s 161570 0 161626 800 6 io_ps[22]
port 222 nsew signal output
rlabel metal2 s 167918 0 167974 800 6 io_ps[23]
port 223 nsew signal output
rlabel metal2 s 174358 0 174414 800 6 io_ps[24]
port 224 nsew signal output
rlabel metal2 s 180798 0 180854 800 6 io_ps[25]
port 225 nsew signal output
rlabel metal2 s 187146 0 187202 800 6 io_ps[26]
port 226 nsew signal output
rlabel metal2 s 193586 0 193642 800 6 io_ps[27]
port 227 nsew signal output
rlabel metal2 s 199934 0 199990 800 6 io_ps[28]
port 228 nsew signal output
rlabel metal2 s 206374 0 206430 800 6 io_ps[29]
port 229 nsew signal output
rlabel metal2 s 33506 0 33562 800 6 io_ps[2]
port 230 nsew signal output
rlabel metal2 s 212722 0 212778 800 6 io_ps[30]
port 231 nsew signal output
rlabel metal2 s 219162 0 219218 800 6 io_ps[31]
port 232 nsew signal output
rlabel metal2 s 39946 0 40002 800 6 io_ps[3]
port 233 nsew signal output
rlabel metal2 s 46386 0 46442 800 6 io_ps[4]
port 234 nsew signal output
rlabel metal2 s 52734 0 52790 800 6 io_ps[5]
port 235 nsew signal output
rlabel metal2 s 59174 0 59230 800 6 io_ps[6]
port 236 nsew signal output
rlabel metal2 s 65522 0 65578 800 6 io_ps[7]
port 237 nsew signal output
rlabel metal2 s 71962 0 72018 800 6 io_ps[8]
port 238 nsew signal output
rlabel metal2 s 78310 0 78366 800 6 io_ps[9]
port 239 nsew signal output
rlabel metal2 s 4710 0 4766 800 6 rst_g
port 240 nsew signal input
rlabel metal2 s 11150 0 11206 800 6 rx
port 241 nsew signal input
rlabel metal2 s 7930 0 7986 800 6 tx
port 242 nsew signal output
rlabel metal3 s 0 4088 800 4208 6 vb_addr0[0]
port 243 nsew signal output
rlabel metal3 s 0 69776 800 69896 6 vb_addr0[10]
port 244 nsew signal output
rlabel metal3 s 0 75896 800 76016 6 vb_addr0[11]
port 245 nsew signal output
rlabel metal3 s 0 82016 800 82136 6 vb_addr0[12]
port 246 nsew signal output
rlabel metal3 s 0 11432 800 11552 6 vb_addr0[1]
port 247 nsew signal output
rlabel metal3 s 0 18776 800 18896 6 vb_addr0[2]
port 248 nsew signal output
rlabel metal3 s 0 25984 800 26104 6 vb_addr0[3]
port 249 nsew signal output
rlabel metal3 s 0 33328 800 33448 6 vb_addr0[4]
port 250 nsew signal output
rlabel metal3 s 0 39448 800 39568 6 vb_addr0[5]
port 251 nsew signal output
rlabel metal3 s 0 45432 800 45552 6 vb_addr0[6]
port 252 nsew signal output
rlabel metal3 s 0 51552 800 51672 6 vb_addr0[7]
port 253 nsew signal output
rlabel metal3 s 0 57672 800 57792 6 vb_addr0[8]
port 254 nsew signal output
rlabel metal3 s 0 63792 800 63912 6 vb_addr0[9]
port 255 nsew signal output
rlabel metal3 s 0 5312 800 5432 6 vb_addr1[0]
port 256 nsew signal output
rlabel metal3 s 0 71000 800 71120 6 vb_addr1[10]
port 257 nsew signal output
rlabel metal3 s 0 77120 800 77240 6 vb_addr1[11]
port 258 nsew signal output
rlabel metal3 s 0 83240 800 83360 6 vb_addr1[12]
port 259 nsew signal output
rlabel metal3 s 0 12656 800 12776 6 vb_addr1[1]
port 260 nsew signal output
rlabel metal3 s 0 20000 800 20120 6 vb_addr1[2]
port 261 nsew signal output
rlabel metal3 s 0 27208 800 27328 6 vb_addr1[3]
port 262 nsew signal output
rlabel metal3 s 0 34552 800 34672 6 vb_addr1[4]
port 263 nsew signal output
rlabel metal3 s 0 40672 800 40792 6 vb_addr1[5]
port 264 nsew signal output
rlabel metal3 s 0 46656 800 46776 6 vb_addr1[6]
port 265 nsew signal output
rlabel metal3 s 0 52776 800 52896 6 vb_addr1[7]
port 266 nsew signal output
rlabel metal3 s 0 58896 800 59016 6 vb_addr1[8]
port 267 nsew signal output
rlabel metal3 s 0 64880 800 65000 6 vb_addr1[9]
port 268 nsew signal output
rlabel metal3 s 0 552 800 672 6 vb_csb0
port 269 nsew signal output
rlabel metal3 s 0 1640 800 1760 6 vb_csb1
port 270 nsew signal output
rlabel metal3 s 0 6536 800 6656 6 vb_din0[0]
port 271 nsew signal output
rlabel metal3 s 0 72224 800 72344 6 vb_din0[10]
port 272 nsew signal output
rlabel metal3 s 0 78344 800 78464 6 vb_din0[11]
port 273 nsew signal output
rlabel metal3 s 0 84464 800 84584 6 vb_din0[12]
port 274 nsew signal output
rlabel metal3 s 0 88000 800 88120 6 vb_din0[13]
port 275 nsew signal output
rlabel metal3 s 0 91672 800 91792 6 vb_din0[14]
port 276 nsew signal output
rlabel metal3 s 0 95344 800 95464 6 vb_din0[15]
port 277 nsew signal output
rlabel metal3 s 0 99016 800 99136 6 vb_din0[16]
port 278 nsew signal output
rlabel metal3 s 0 102688 800 102808 6 vb_din0[17]
port 279 nsew signal output
rlabel metal3 s 0 106360 800 106480 6 vb_din0[18]
port 280 nsew signal output
rlabel metal3 s 0 109896 800 110016 6 vb_din0[19]
port 281 nsew signal output
rlabel metal3 s 0 13880 800 14000 6 vb_din0[1]
port 282 nsew signal output
rlabel metal3 s 0 113568 800 113688 6 vb_din0[20]
port 283 nsew signal output
rlabel metal3 s 0 117240 800 117360 6 vb_din0[21]
port 284 nsew signal output
rlabel metal3 s 0 120912 800 121032 6 vb_din0[22]
port 285 nsew signal output
rlabel metal3 s 0 124584 800 124704 6 vb_din0[23]
port 286 nsew signal output
rlabel metal3 s 0 128120 800 128240 6 vb_din0[24]
port 287 nsew signal output
rlabel metal3 s 0 131792 800 131912 6 vb_din0[25]
port 288 nsew signal output
rlabel metal3 s 0 135464 800 135584 6 vb_din0[26]
port 289 nsew signal output
rlabel metal3 s 0 139136 800 139256 6 vb_din0[27]
port 290 nsew signal output
rlabel metal3 s 0 142808 800 142928 6 vb_din0[28]
port 291 nsew signal output
rlabel metal3 s 0 146480 800 146600 6 vb_din0[29]
port 292 nsew signal output
rlabel metal3 s 0 21224 800 21344 6 vb_din0[2]
port 293 nsew signal output
rlabel metal3 s 0 150016 800 150136 6 vb_din0[30]
port 294 nsew signal output
rlabel metal3 s 0 153688 800 153808 6 vb_din0[31]
port 295 nsew signal output
rlabel metal3 s 0 28432 800 28552 6 vb_din0[3]
port 296 nsew signal output
rlabel metal3 s 0 35776 800 35896 6 vb_din0[4]
port 297 nsew signal output
rlabel metal3 s 0 41896 800 42016 6 vb_din0[5]
port 298 nsew signal output
rlabel metal3 s 0 47880 800 48000 6 vb_din0[6]
port 299 nsew signal output
rlabel metal3 s 0 54000 800 54120 6 vb_din0[7]
port 300 nsew signal output
rlabel metal3 s 0 60120 800 60240 6 vb_din0[8]
port 301 nsew signal output
rlabel metal3 s 0 66104 800 66224 6 vb_din0[9]
port 302 nsew signal output
rlabel metal3 s 0 7760 800 7880 6 vb_dout0[0]
port 303 nsew signal input
rlabel metal3 s 0 73448 800 73568 6 vb_dout0[10]
port 304 nsew signal input
rlabel metal3 s 0 79568 800 79688 6 vb_dout0[11]
port 305 nsew signal input
rlabel metal3 s 0 85552 800 85672 6 vb_dout0[12]
port 306 nsew signal input
rlabel metal3 s 0 89224 800 89344 6 vb_dout0[13]
port 307 nsew signal input
rlabel metal3 s 0 92896 800 93016 6 vb_dout0[14]
port 308 nsew signal input
rlabel metal3 s 0 96568 800 96688 6 vb_dout0[15]
port 309 nsew signal input
rlabel metal3 s 0 100240 800 100360 6 vb_dout0[16]
port 310 nsew signal input
rlabel metal3 s 0 103912 800 104032 6 vb_dout0[17]
port 311 nsew signal input
rlabel metal3 s 0 107448 800 107568 6 vb_dout0[18]
port 312 nsew signal input
rlabel metal3 s 0 111120 800 111240 6 vb_dout0[19]
port 313 nsew signal input
rlabel metal3 s 0 15104 800 15224 6 vb_dout0[1]
port 314 nsew signal input
rlabel metal3 s 0 114792 800 114912 6 vb_dout0[20]
port 315 nsew signal input
rlabel metal3 s 0 118464 800 118584 6 vb_dout0[21]
port 316 nsew signal input
rlabel metal3 s 0 122136 800 122256 6 vb_dout0[22]
port 317 nsew signal input
rlabel metal3 s 0 125808 800 125928 6 vb_dout0[23]
port 318 nsew signal input
rlabel metal3 s 0 129344 800 129464 6 vb_dout0[24]
port 319 nsew signal input
rlabel metal3 s 0 133016 800 133136 6 vb_dout0[25]
port 320 nsew signal input
rlabel metal3 s 0 136688 800 136808 6 vb_dout0[26]
port 321 nsew signal input
rlabel metal3 s 0 140360 800 140480 6 vb_dout0[27]
port 322 nsew signal input
rlabel metal3 s 0 144032 800 144152 6 vb_dout0[28]
port 323 nsew signal input
rlabel metal3 s 0 147704 800 147824 6 vb_dout0[29]
port 324 nsew signal input
rlabel metal3 s 0 22312 800 22432 6 vb_dout0[2]
port 325 nsew signal input
rlabel metal3 s 0 151240 800 151360 6 vb_dout0[30]
port 326 nsew signal input
rlabel metal3 s 0 154912 800 155032 6 vb_dout0[31]
port 327 nsew signal input
rlabel metal3 s 0 29656 800 29776 6 vb_dout0[3]
port 328 nsew signal input
rlabel metal3 s 0 37000 800 37120 6 vb_dout0[4]
port 329 nsew signal input
rlabel metal3 s 0 42984 800 43104 6 vb_dout0[5]
port 330 nsew signal input
rlabel metal3 s 0 49104 800 49224 6 vb_dout0[6]
port 331 nsew signal input
rlabel metal3 s 0 55224 800 55344 6 vb_dout0[7]
port 332 nsew signal input
rlabel metal3 s 0 61344 800 61464 6 vb_dout0[8]
port 333 nsew signal input
rlabel metal3 s 0 67328 800 67448 6 vb_dout0[9]
port 334 nsew signal input
rlabel metal3 s 0 8984 800 9104 6 vb_dout1[0]
port 335 nsew signal input
rlabel metal3 s 0 74672 800 74792 6 vb_dout1[10]
port 336 nsew signal input
rlabel metal3 s 0 80792 800 80912 6 vb_dout1[11]
port 337 nsew signal input
rlabel metal3 s 0 86776 800 86896 6 vb_dout1[12]
port 338 nsew signal input
rlabel metal3 s 0 90448 800 90568 6 vb_dout1[13]
port 339 nsew signal input
rlabel metal3 s 0 94120 800 94240 6 vb_dout1[14]
port 340 nsew signal input
rlabel metal3 s 0 97792 800 97912 6 vb_dout1[15]
port 341 nsew signal input
rlabel metal3 s 0 101464 800 101584 6 vb_dout1[16]
port 342 nsew signal input
rlabel metal3 s 0 105136 800 105256 6 vb_dout1[17]
port 343 nsew signal input
rlabel metal3 s 0 108672 800 108792 6 vb_dout1[18]
port 344 nsew signal input
rlabel metal3 s 0 112344 800 112464 6 vb_dout1[19]
port 345 nsew signal input
rlabel metal3 s 0 16328 800 16448 6 vb_dout1[1]
port 346 nsew signal input
rlabel metal3 s 0 116016 800 116136 6 vb_dout1[20]
port 347 nsew signal input
rlabel metal3 s 0 119688 800 119808 6 vb_dout1[21]
port 348 nsew signal input
rlabel metal3 s 0 123360 800 123480 6 vb_dout1[22]
port 349 nsew signal input
rlabel metal3 s 0 127032 800 127152 6 vb_dout1[23]
port 350 nsew signal input
rlabel metal3 s 0 130568 800 130688 6 vb_dout1[24]
port 351 nsew signal input
rlabel metal3 s 0 134240 800 134360 6 vb_dout1[25]
port 352 nsew signal input
rlabel metal3 s 0 137912 800 138032 6 vb_dout1[26]
port 353 nsew signal input
rlabel metal3 s 0 141584 800 141704 6 vb_dout1[27]
port 354 nsew signal input
rlabel metal3 s 0 145256 800 145376 6 vb_dout1[28]
port 355 nsew signal input
rlabel metal3 s 0 148792 800 148912 6 vb_dout1[29]
port 356 nsew signal input
rlabel metal3 s 0 23536 800 23656 6 vb_dout1[2]
port 357 nsew signal input
rlabel metal3 s 0 152464 800 152584 6 vb_dout1[30]
port 358 nsew signal input
rlabel metal3 s 0 156136 800 156256 6 vb_dout1[31]
port 359 nsew signal input
rlabel metal3 s 0 30880 800 31000 6 vb_dout1[3]
port 360 nsew signal input
rlabel metal3 s 0 38224 800 38344 6 vb_dout1[4]
port 361 nsew signal input
rlabel metal3 s 0 44208 800 44328 6 vb_dout1[5]
port 362 nsew signal input
rlabel metal3 s 0 50328 800 50448 6 vb_dout1[6]
port 363 nsew signal input
rlabel metal3 s 0 56448 800 56568 6 vb_dout1[7]
port 364 nsew signal input
rlabel metal3 s 0 62568 800 62688 6 vb_dout1[8]
port 365 nsew signal input
rlabel metal3 s 0 68552 800 68672 6 vb_dout1[9]
port 366 nsew signal input
rlabel metal3 s 0 2864 800 2984 6 vb_web0
port 367 nsew signal output
rlabel metal3 s 0 10208 800 10328 6 vb_wmask0[0]
port 368 nsew signal output
rlabel metal3 s 0 17552 800 17672 6 vb_wmask0[1]
port 369 nsew signal output
rlabel metal3 s 0 24760 800 24880 6 vb_wmask0[2]
port 370 nsew signal output
rlabel metal3 s 0 32104 800 32224 6 vb_wmask0[3]
port 371 nsew signal output
rlabel metal4 s 4208 2128 4528 357456 6 vccd1
port 372 nsew power input
rlabel metal4 s 34928 2128 35248 357456 6 vccd1
port 372 nsew power input
rlabel metal4 s 65648 2128 65968 357456 6 vccd1
port 372 nsew power input
rlabel metal4 s 96368 2128 96688 357456 6 vccd1
port 372 nsew power input
rlabel metal4 s 127088 2128 127408 357456 6 vccd1
port 372 nsew power input
rlabel metal4 s 157808 2128 158128 357456 6 vccd1
port 372 nsew power input
rlabel metal4 s 188528 2128 188848 357456 6 vccd1
port 372 nsew power input
rlabel metal4 s 219248 2128 219568 357456 6 vccd1
port 372 nsew power input
rlabel metal4 s 19568 2128 19888 357456 6 vssd1
port 373 nsew ground input
rlabel metal4 s 50288 2128 50608 357456 6 vssd1
port 373 nsew ground input
rlabel metal4 s 81008 2128 81328 357456 6 vssd1
port 373 nsew ground input
rlabel metal4 s 111728 2128 112048 357456 6 vssd1
port 373 nsew ground input
rlabel metal4 s 142448 2128 142768 357456 6 vssd1
port 373 nsew ground input
rlabel metal4 s 173168 2128 173488 357456 6 vssd1
port 373 nsew ground input
rlabel metal4 s 203888 2128 204208 357456 6 vssd1
port 373 nsew ground input
rlabel metal4 s 234608 2128 234928 357456 6 vssd1
port 373 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 240000 360000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 75858108
string GDS_FILE /home/kasirga/c0_hayyan/GL_GECTI/caravel_user_project/openlane/c0_system/runs/c0_system/results/finishing/c0_system.magic.gds
string GDS_START 1677124
<< end >>


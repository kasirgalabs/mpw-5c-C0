VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO c0_system
  CLASS BLOCK ;
  FOREIGN c0_system ;
  ORIGIN 0.000 0.000 ;
  SIZE 1500.000 BY 1500.000 ;
  PIN bb_addr0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 670.520 4.000 671.120 ;
    END
  END bb_addr0[0]
  PIN bb_addr0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 944.560 4.000 945.160 ;
    END
  END bb_addr0[10]
  PIN bb_addr0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 969.720 4.000 970.320 ;
    END
  END bb_addr0[11]
  PIN bb_addr0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 994.880 4.000 995.480 ;
    END
  END bb_addr0[12]
  PIN bb_addr0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1020.040 4.000 1020.640 ;
    END
  END bb_addr0[13]
  PIN bb_addr0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1045.880 4.000 1046.480 ;
    END
  END bb_addr0[14]
  PIN bb_addr0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1071.040 4.000 1071.640 ;
    END
  END bb_addr0[15]
  PIN bb_addr0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1096.200 4.000 1096.800 ;
    END
  END bb_addr0[16]
  PIN bb_addr0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1122.040 4.000 1122.640 ;
    END
  END bb_addr0[17]
  PIN bb_addr0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1147.200 4.000 1147.800 ;
    END
  END bb_addr0[18]
  PIN bb_addr0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1172.360 4.000 1172.960 ;
    END
  END bb_addr0[19]
  PIN bb_addr0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 701.120 4.000 701.720 ;
    END
  END bb_addr0[1]
  PIN bb_addr0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1197.520 4.000 1198.120 ;
    END
  END bb_addr0[20]
  PIN bb_addr0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1223.360 4.000 1223.960 ;
    END
  END bb_addr0[21]
  PIN bb_addr0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1248.520 4.000 1249.120 ;
    END
  END bb_addr0[22]
  PIN bb_addr0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1273.680 4.000 1274.280 ;
    END
  END bb_addr0[23]
  PIN bb_addr0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1298.840 4.000 1299.440 ;
    END
  END bb_addr0[24]
  PIN bb_addr0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1324.680 4.000 1325.280 ;
    END
  END bb_addr0[25]
  PIN bb_addr0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1349.840 4.000 1350.440 ;
    END
  END bb_addr0[26]
  PIN bb_addr0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1375.000 4.000 1375.600 ;
    END
  END bb_addr0[27]
  PIN bb_addr0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1400.160 4.000 1400.760 ;
    END
  END bb_addr0[28]
  PIN bb_addr0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1426.000 4.000 1426.600 ;
    END
  END bb_addr0[29]
  PIN bb_addr0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 731.720 4.000 732.320 ;
    END
  END bb_addr0[2]
  PIN bb_addr0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1451.160 4.000 1451.760 ;
    END
  END bb_addr0[30]
  PIN bb_addr0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1476.320 4.000 1476.920 ;
    END
  END bb_addr0[31]
  PIN bb_addr0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 761.640 4.000 762.240 ;
    END
  END bb_addr0[3]
  PIN bb_addr0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 792.240 4.000 792.840 ;
    END
  END bb_addr0[4]
  PIN bb_addr0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 817.400 4.000 818.000 ;
    END
  END bb_addr0[5]
  PIN bb_addr0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 843.240 4.000 843.840 ;
    END
  END bb_addr0[6]
  PIN bb_addr0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 868.400 4.000 869.000 ;
    END
  END bb_addr0[7]
  PIN bb_addr0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 893.560 4.000 894.160 ;
    END
  END bb_addr0[8]
  PIN bb_addr0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 918.720 4.000 919.320 ;
    END
  END bb_addr0[9]
  PIN bb_addr1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 675.960 4.000 676.560 ;
    END
  END bb_addr1[0]
  PIN bb_addr1[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 949.320 4.000 949.920 ;
    END
  END bb_addr1[10]
  PIN bb_addr1[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 974.480 4.000 975.080 ;
    END
  END bb_addr1[11]
  PIN bb_addr1[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1000.320 4.000 1000.920 ;
    END
  END bb_addr1[12]
  PIN bb_addr1[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1025.480 4.000 1026.080 ;
    END
  END bb_addr1[13]
  PIN bb_addr1[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1050.640 4.000 1051.240 ;
    END
  END bb_addr1[14]
  PIN bb_addr1[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1075.800 4.000 1076.400 ;
    END
  END bb_addr1[15]
  PIN bb_addr1[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1101.640 4.000 1102.240 ;
    END
  END bb_addr1[16]
  PIN bb_addr1[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1126.800 4.000 1127.400 ;
    END
  END bb_addr1[17]
  PIN bb_addr1[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1151.960 4.000 1152.560 ;
    END
  END bb_addr1[18]
  PIN bb_addr1[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1177.800 4.000 1178.400 ;
    END
  END bb_addr1[19]
  PIN bb_addr1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 705.880 4.000 706.480 ;
    END
  END bb_addr1[1]
  PIN bb_addr1[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1202.960 4.000 1203.560 ;
    END
  END bb_addr1[20]
  PIN bb_addr1[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1228.120 4.000 1228.720 ;
    END
  END bb_addr1[21]
  PIN bb_addr1[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1253.280 4.000 1253.880 ;
    END
  END bb_addr1[22]
  PIN bb_addr1[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1279.120 4.000 1279.720 ;
    END
  END bb_addr1[23]
  PIN bb_addr1[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1304.280 4.000 1304.880 ;
    END
  END bb_addr1[24]
  PIN bb_addr1[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1329.440 4.000 1330.040 ;
    END
  END bb_addr1[25]
  PIN bb_addr1[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1354.600 4.000 1355.200 ;
    END
  END bb_addr1[26]
  PIN bb_addr1[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1380.440 4.000 1381.040 ;
    END
  END bb_addr1[27]
  PIN bb_addr1[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1405.600 4.000 1406.200 ;
    END
  END bb_addr1[28]
  PIN bb_addr1[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1430.760 4.000 1431.360 ;
    END
  END bb_addr1[29]
  PIN bb_addr1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 736.480 4.000 737.080 ;
    END
  END bb_addr1[2]
  PIN bb_addr1[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1455.920 4.000 1456.520 ;
    END
  END bb_addr1[30]
  PIN bb_addr1[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1481.760 4.000 1482.360 ;
    END
  END bb_addr1[31]
  PIN bb_addr1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 767.080 4.000 767.680 ;
    END
  END bb_addr1[3]
  PIN bb_addr1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 797.680 4.000 798.280 ;
    END
  END bb_addr1[4]
  PIN bb_addr1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 822.840 4.000 823.440 ;
    END
  END bb_addr1[5]
  PIN bb_addr1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 848.000 4.000 848.600 ;
    END
  END bb_addr1[6]
  PIN bb_addr1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 873.160 4.000 873.760 ;
    END
  END bb_addr1[7]
  PIN bb_addr1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 899.000 4.000 899.600 ;
    END
  END bb_addr1[8]
  PIN bb_addr1[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 924.160 4.000 924.760 ;
    END
  END bb_addr1[9]
  PIN bb_csb0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 655.560 4.000 656.160 ;
    END
  END bb_csb0
  PIN bb_csb1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 660.320 4.000 660.920 ;
    END
  END bb_csb1
  PIN bb_din0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 680.720 4.000 681.320 ;
    END
  END bb_din0[0]
  PIN bb_din0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 954.760 4.000 955.360 ;
    END
  END bb_din0[10]
  PIN bb_din0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 979.920 4.000 980.520 ;
    END
  END bb_din0[11]
  PIN bb_din0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1005.080 4.000 1005.680 ;
    END
  END bb_din0[12]
  PIN bb_din0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1030.240 4.000 1030.840 ;
    END
  END bb_din0[13]
  PIN bb_din0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1056.080 4.000 1056.680 ;
    END
  END bb_din0[14]
  PIN bb_din0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1081.240 4.000 1081.840 ;
    END
  END bb_din0[15]
  PIN bb_din0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1106.400 4.000 1107.000 ;
    END
  END bb_din0[16]
  PIN bb_din0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1131.560 4.000 1132.160 ;
    END
  END bb_din0[17]
  PIN bb_din0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1157.400 4.000 1158.000 ;
    END
  END bb_din0[18]
  PIN bb_din0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1182.560 4.000 1183.160 ;
    END
  END bb_din0[19]
  PIN bb_din0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 711.320 4.000 711.920 ;
    END
  END bb_din0[1]
  PIN bb_din0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1207.720 4.000 1208.320 ;
    END
  END bb_din0[20]
  PIN bb_din0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1233.560 4.000 1234.160 ;
    END
  END bb_din0[21]
  PIN bb_din0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1258.720 4.000 1259.320 ;
    END
  END bb_din0[22]
  PIN bb_din0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1283.880 4.000 1284.480 ;
    END
  END bb_din0[23]
  PIN bb_din0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1309.040 4.000 1309.640 ;
    END
  END bb_din0[24]
  PIN bb_din0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1334.880 4.000 1335.480 ;
    END
  END bb_din0[25]
  PIN bb_din0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1360.040 4.000 1360.640 ;
    END
  END bb_din0[26]
  PIN bb_din0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1385.200 4.000 1385.800 ;
    END
  END bb_din0[27]
  PIN bb_din0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1410.360 4.000 1410.960 ;
    END
  END bb_din0[28]
  PIN bb_din0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1436.200 4.000 1436.800 ;
    END
  END bb_din0[29]
  PIN bb_din0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 741.920 4.000 742.520 ;
    END
  END bb_din0[2]
  PIN bb_din0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1461.360 4.000 1461.960 ;
    END
  END bb_din0[30]
  PIN bb_din0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1486.520 4.000 1487.120 ;
    END
  END bb_din0[31]
  PIN bb_din0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 771.840 4.000 772.440 ;
    END
  END bb_din0[3]
  PIN bb_din0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 802.440 4.000 803.040 ;
    END
  END bb_din0[4]
  PIN bb_din0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 827.600 4.000 828.200 ;
    END
  END bb_din0[5]
  PIN bb_din0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 853.440 4.000 854.040 ;
    END
  END bb_din0[6]
  PIN bb_din0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 878.600 4.000 879.200 ;
    END
  END bb_din0[7]
  PIN bb_din0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 903.760 4.000 904.360 ;
    END
  END bb_din0[8]
  PIN bb_din0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 928.920 4.000 929.520 ;
    END
  END bb_din0[9]
  PIN bb_dout0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 686.160 4.000 686.760 ;
    END
  END bb_dout0[0]
  PIN bb_dout0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 959.520 4.000 960.120 ;
    END
  END bb_dout0[10]
  PIN bb_dout0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 984.680 4.000 985.280 ;
    END
  END bb_dout0[11]
  PIN bb_dout0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1010.520 4.000 1011.120 ;
    END
  END bb_dout0[12]
  PIN bb_dout0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1035.680 4.000 1036.280 ;
    END
  END bb_dout0[13]
  PIN bb_dout0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1060.840 4.000 1061.440 ;
    END
  END bb_dout0[14]
  PIN bb_dout0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1086.000 4.000 1086.600 ;
    END
  END bb_dout0[15]
  PIN bb_dout0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1111.840 4.000 1112.440 ;
    END
  END bb_dout0[16]
  PIN bb_dout0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1137.000 4.000 1137.600 ;
    END
  END bb_dout0[17]
  PIN bb_dout0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1162.160 4.000 1162.760 ;
    END
  END bb_dout0[18]
  PIN bb_dout0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1187.320 4.000 1187.920 ;
    END
  END bb_dout0[19]
  PIN bb_dout0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 716.080 4.000 716.680 ;
    END
  END bb_dout0[1]
  PIN bb_dout0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1213.160 4.000 1213.760 ;
    END
  END bb_dout0[20]
  PIN bb_dout0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1238.320 4.000 1238.920 ;
    END
  END bb_dout0[21]
  PIN bb_dout0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1263.480 4.000 1264.080 ;
    END
  END bb_dout0[22]
  PIN bb_dout0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1288.640 4.000 1289.240 ;
    END
  END bb_dout0[23]
  PIN bb_dout0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1314.480 4.000 1315.080 ;
    END
  END bb_dout0[24]
  PIN bb_dout0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1339.640 4.000 1340.240 ;
    END
  END bb_dout0[25]
  PIN bb_dout0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1364.800 4.000 1365.400 ;
    END
  END bb_dout0[26]
  PIN bb_dout0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1390.640 4.000 1391.240 ;
    END
  END bb_dout0[27]
  PIN bb_dout0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1415.800 4.000 1416.400 ;
    END
  END bb_dout0[28]
  PIN bb_dout0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1440.960 4.000 1441.560 ;
    END
  END bb_dout0[29]
  PIN bb_dout0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 746.680 4.000 747.280 ;
    END
  END bb_dout0[2]
  PIN bb_dout0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1466.120 4.000 1466.720 ;
    END
  END bb_dout0[30]
  PIN bb_dout0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1491.960 4.000 1492.560 ;
    END
  END bb_dout0[31]
  PIN bb_dout0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 777.280 4.000 777.880 ;
    END
  END bb_dout0[3]
  PIN bb_dout0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 807.200 4.000 807.800 ;
    END
  END bb_dout0[4]
  PIN bb_dout0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 833.040 4.000 833.640 ;
    END
  END bb_dout0[5]
  PIN bb_dout0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 858.200 4.000 858.800 ;
    END
  END bb_dout0[6]
  PIN bb_dout0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 883.360 4.000 883.960 ;
    END
  END bb_dout0[7]
  PIN bb_dout0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 909.200 4.000 909.800 ;
    END
  END bb_dout0[8]
  PIN bb_dout0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 934.360 4.000 934.960 ;
    END
  END bb_dout0[9]
  PIN bb_dout1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 690.920 4.000 691.520 ;
    END
  END bb_dout1[0]
  PIN bb_dout1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 964.960 4.000 965.560 ;
    END
  END bb_dout1[10]
  PIN bb_dout1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 990.120 4.000 990.720 ;
    END
  END bb_dout1[11]
  PIN bb_dout1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1015.280 4.000 1015.880 ;
    END
  END bb_dout1[12]
  PIN bb_dout1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1040.440 4.000 1041.040 ;
    END
  END bb_dout1[13]
  PIN bb_dout1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1066.280 4.000 1066.880 ;
    END
  END bb_dout1[14]
  PIN bb_dout1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1091.440 4.000 1092.040 ;
    END
  END bb_dout1[15]
  PIN bb_dout1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1116.600 4.000 1117.200 ;
    END
  END bb_dout1[16]
  PIN bb_dout1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1141.760 4.000 1142.360 ;
    END
  END bb_dout1[17]
  PIN bb_dout1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1167.600 4.000 1168.200 ;
    END
  END bb_dout1[18]
  PIN bb_dout1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1192.760 4.000 1193.360 ;
    END
  END bb_dout1[19]
  PIN bb_dout1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 721.520 4.000 722.120 ;
    END
  END bb_dout1[1]
  PIN bb_dout1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1217.920 4.000 1218.520 ;
    END
  END bb_dout1[20]
  PIN bb_dout1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1243.080 4.000 1243.680 ;
    END
  END bb_dout1[21]
  PIN bb_dout1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1268.920 4.000 1269.520 ;
    END
  END bb_dout1[22]
  PIN bb_dout1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1294.080 4.000 1294.680 ;
    END
  END bb_dout1[23]
  PIN bb_dout1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1319.240 4.000 1319.840 ;
    END
  END bb_dout1[24]
  PIN bb_dout1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1344.400 4.000 1345.000 ;
    END
  END bb_dout1[25]
  PIN bb_dout1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1370.240 4.000 1370.840 ;
    END
  END bb_dout1[26]
  PIN bb_dout1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1395.400 4.000 1396.000 ;
    END
  END bb_dout1[27]
  PIN bb_dout1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1420.560 4.000 1421.160 ;
    END
  END bb_dout1[28]
  PIN bb_dout1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1446.400 4.000 1447.000 ;
    END
  END bb_dout1[29]
  PIN bb_dout1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 752.120 4.000 752.720 ;
    END
  END bb_dout1[2]
  PIN bb_dout1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1471.560 4.000 1472.160 ;
    END
  END bb_dout1[30]
  PIN bb_dout1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1496.720 4.000 1497.320 ;
    END
  END bb_dout1[31]
  PIN bb_dout1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 782.040 4.000 782.640 ;
    END
  END bb_dout1[3]
  PIN bb_dout1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 812.640 4.000 813.240 ;
    END
  END bb_dout1[4]
  PIN bb_dout1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 837.800 4.000 838.400 ;
    END
  END bb_dout1[5]
  PIN bb_dout1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 862.960 4.000 863.560 ;
    END
  END bb_dout1[6]
  PIN bb_dout1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 888.800 4.000 889.400 ;
    END
  END bb_dout1[7]
  PIN bb_dout1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 913.960 4.000 914.560 ;
    END
  END bb_dout1[8]
  PIN bb_dout1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 939.120 4.000 939.720 ;
    END
  END bb_dout1[9]
  PIN bb_web0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 665.760 4.000 666.360 ;
    END
  END bb_web0
  PIN bb_wmask0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 696.360 4.000 696.960 ;
    END
  END bb_wmask0[0]
  PIN bb_wmask0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 726.280 4.000 726.880 ;
    END
  END bb_wmask0[1]
  PIN bb_wmask0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 756.880 4.000 757.480 ;
    END
  END bb_wmask0[2]
  PIN bb_wmask0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 787.480 4.000 788.080 ;
    END
  END bb_wmask0[3]
  PIN clk_g
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 0.000 10.030 4.000 ;
    END
  END clk_g
  PIN io_gecerli
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.330 0.000 89.610 4.000 ;
    END
  END io_gecerli
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 4.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 509.770 0.000 510.050 4.000 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 549.330 0.000 549.610 4.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 589.350 0.000 589.630 4.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 629.370 0.000 629.650 4.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 669.390 0.000 669.670 4.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 709.410 0.000 709.690 4.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 749.430 0.000 749.710 4.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 789.450 0.000 789.730 4.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 829.470 0.000 829.750 4.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 869.490 0.000 869.770 4.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.590 0.000 149.870 4.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 909.510 0.000 909.790 4.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 949.530 0.000 949.810 4.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 989.550 0.000 989.830 4.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1029.570 0.000 1029.850 4.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1069.590 0.000 1069.870 4.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1109.610 0.000 1109.890 4.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1149.630 0.000 1149.910 4.000 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1189.650 0.000 1189.930 4.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1229.670 0.000 1229.950 4.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1269.690 0.000 1269.970 4.000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.610 0.000 189.890 4.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1309.710 0.000 1309.990 4.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1349.730 0.000 1350.010 4.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1389.750 0.000 1390.030 4.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1409.530 0.000 1409.810 4.000 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1429.770 0.000 1430.050 4.000 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1449.550 0.000 1449.830 4.000 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1469.790 0.000 1470.070 4.000 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1489.570 0.000 1489.850 4.000 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.630 0.000 229.910 4.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.650 0.000 269.930 4.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.670 0.000 309.950 4.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 349.690 0.000 349.970 4.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.710 0.000 389.990 4.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 429.730 0.000 430.010 4.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 469.750 0.000 470.030 4.000 ;
    END
  END io_oeb[9]
  PIN io_ps[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.350 0.000 129.630 4.000 ;
    END
  END io_ps[0]
  PIN io_ps[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 529.550 0.000 529.830 4.000 ;
    END
  END io_ps[10]
  PIN io_ps[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 569.570 0.000 569.850 4.000 ;
    END
  END io_ps[11]
  PIN io_ps[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 609.590 0.000 609.870 4.000 ;
    END
  END io_ps[12]
  PIN io_ps[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 649.610 0.000 649.890 4.000 ;
    END
  END io_ps[13]
  PIN io_ps[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 689.630 0.000 689.910 4.000 ;
    END
  END io_ps[14]
  PIN io_ps[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 729.650 0.000 729.930 4.000 ;
    END
  END io_ps[15]
  PIN io_ps[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 769.670 0.000 769.950 4.000 ;
    END
  END io_ps[16]
  PIN io_ps[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 809.690 0.000 809.970 4.000 ;
    END
  END io_ps[17]
  PIN io_ps[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 849.710 0.000 849.990 4.000 ;
    END
  END io_ps[18]
  PIN io_ps[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 889.730 0.000 890.010 4.000 ;
    END
  END io_ps[19]
  PIN io_ps[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.370 0.000 169.650 4.000 ;
    END
  END io_ps[1]
  PIN io_ps[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 929.750 0.000 930.030 4.000 ;
    END
  END io_ps[20]
  PIN io_ps[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 969.770 0.000 970.050 4.000 ;
    END
  END io_ps[21]
  PIN io_ps[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1009.790 0.000 1010.070 4.000 ;
    END
  END io_ps[22]
  PIN io_ps[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1049.350 0.000 1049.630 4.000 ;
    END
  END io_ps[23]
  PIN io_ps[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1089.370 0.000 1089.650 4.000 ;
    END
  END io_ps[24]
  PIN io_ps[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1129.390 0.000 1129.670 4.000 ;
    END
  END io_ps[25]
  PIN io_ps[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1169.410 0.000 1169.690 4.000 ;
    END
  END io_ps[26]
  PIN io_ps[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1209.430 0.000 1209.710 4.000 ;
    END
  END io_ps[27]
  PIN io_ps[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1249.450 0.000 1249.730 4.000 ;
    END
  END io_ps[28]
  PIN io_ps[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1289.470 0.000 1289.750 4.000 ;
    END
  END io_ps[29]
  PIN io_ps[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.390 0.000 209.670 4.000 ;
    END
  END io_ps[2]
  PIN io_ps[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1329.490 0.000 1329.770 4.000 ;
    END
  END io_ps[30]
  PIN io_ps[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1369.510 0.000 1369.790 4.000 ;
    END
  END io_ps[31]
  PIN io_ps[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.410 0.000 249.690 4.000 ;
    END
  END io_ps[3]
  PIN io_ps[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.430 0.000 289.710 4.000 ;
    END
  END io_ps[4]
  PIN io_ps[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 329.450 0.000 329.730 4.000 ;
    END
  END io_ps[5]
  PIN io_ps[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.470 0.000 369.750 4.000 ;
    END
  END io_ps[6]
  PIN io_ps[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.490 0.000 409.770 4.000 ;
    END
  END io_ps[7]
  PIN io_ps[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.510 0.000 449.790 4.000 ;
    END
  END io_ps[8]
  PIN io_ps[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.530 0.000 489.810 4.000 ;
    END
  END io_ps[9]
  PIN rst_g
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.530 0.000 29.810 4.000 ;
    END
  END rst_g
  PIN rx
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.550 0.000 69.830 4.000 ;
    END
  END rx
  PIN tx
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.310 0.000 49.590 4.000 ;
    END
  END tx
  PIN vb_addr0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 4.000 17.640 ;
    END
  END vb_addr0[0]
  PIN vb_addr0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 290.400 4.000 291.000 ;
    END
  END vb_addr0[10]
  PIN vb_addr0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 316.240 4.000 316.840 ;
    END
  END vb_addr0[11]
  PIN vb_addr0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 341.400 4.000 342.000 ;
    END
  END vb_addr0[12]
  PIN vb_addr0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END vb_addr0[1]
  PIN vb_addr0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 77.560 4.000 78.160 ;
    END
  END vb_addr0[2]
  PIN vb_addr0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.160 4.000 108.760 ;
    END
  END vb_addr0[3]
  PIN vb_addr0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 138.760 4.000 139.360 ;
    END
  END vb_addr0[4]
  PIN vb_addr0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.920 4.000 164.520 ;
    END
  END vb_addr0[5]
  PIN vb_addr0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 189.080 4.000 189.680 ;
    END
  END vb_addr0[6]
  PIN vb_addr0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.920 4.000 215.520 ;
    END
  END vb_addr0[7]
  PIN vb_addr0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 240.080 4.000 240.680 ;
    END
  END vb_addr0[8]
  PIN vb_addr0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 265.240 4.000 265.840 ;
    END
  END vb_addr0[9]
  PIN vb_addr1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.800 4.000 22.400 ;
    END
  END vb_addr1[0]
  PIN vb_addr1[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 295.840 4.000 296.440 ;
    END
  END vb_addr1[10]
  PIN vb_addr1[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 321.000 4.000 321.600 ;
    END
  END vb_addr1[11]
  PIN vb_addr1[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 346.160 4.000 346.760 ;
    END
  END vb_addr1[12]
  PIN vb_addr1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 52.400 4.000 53.000 ;
    END
  END vb_addr1[1]
  PIN vb_addr1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.000 4.000 83.600 ;
    END
  END vb_addr1[2]
  PIN vb_addr1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.920 4.000 113.520 ;
    END
  END vb_addr1[3]
  PIN vb_addr1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 143.520 4.000 144.120 ;
    END
  END vb_addr1[4]
  PIN vb_addr1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.680 4.000 169.280 ;
    END
  END vb_addr1[5]
  PIN vb_addr1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 194.520 4.000 195.120 ;
    END
  END vb_addr1[6]
  PIN vb_addr1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 219.680 4.000 220.280 ;
    END
  END vb_addr1[7]
  PIN vb_addr1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 244.840 4.000 245.440 ;
    END
  END vb_addr1[8]
  PIN vb_addr1[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 270.000 4.000 270.600 ;
    END
  END vb_addr1[9]
  PIN vb_csb0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.080 4.000 2.680 ;
    END
  END vb_csb0
  PIN vb_csb1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END vb_csb1
  PIN vb_din0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END vb_din0[0]
  PIN vb_din0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 300.600 4.000 301.200 ;
    END
  END vb_din0[10]
  PIN vb_din0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 325.760 4.000 326.360 ;
    END
  END vb_din0[11]
  PIN vb_din0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 351.600 4.000 352.200 ;
    END
  END vb_din0[12]
  PIN vb_din0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 366.560 4.000 367.160 ;
    END
  END vb_din0[13]
  PIN vb_din0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 381.520 4.000 382.120 ;
    END
  END vb_din0[14]
  PIN vb_din0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 397.160 4.000 397.760 ;
    END
  END vb_din0[15]
  PIN vb_din0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 412.120 4.000 412.720 ;
    END
  END vb_din0[16]
  PIN vb_din0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 427.760 4.000 428.360 ;
    END
  END vb_din0[17]
  PIN vb_din0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 442.720 4.000 443.320 ;
    END
  END vb_din0[18]
  PIN vb_din0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 457.680 4.000 458.280 ;
    END
  END vb_din0[19]
  PIN vb_din0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.160 4.000 57.760 ;
    END
  END vb_din0[1]
  PIN vb_din0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 473.320 4.000 473.920 ;
    END
  END vb_din0[20]
  PIN vb_din0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 488.280 4.000 488.880 ;
    END
  END vb_din0[21]
  PIN vb_din0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 503.240 4.000 503.840 ;
    END
  END vb_din0[22]
  PIN vb_din0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 518.880 4.000 519.480 ;
    END
  END vb_din0[23]
  PIN vb_din0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 533.840 4.000 534.440 ;
    END
  END vb_din0[24]
  PIN vb_din0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 548.800 4.000 549.400 ;
    END
  END vb_din0[25]
  PIN vb_din0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 564.440 4.000 565.040 ;
    END
  END vb_din0[26]
  PIN vb_din0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 579.400 4.000 580.000 ;
    END
  END vb_din0[27]
  PIN vb_din0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 594.360 4.000 594.960 ;
    END
  END vb_din0[28]
  PIN vb_din0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 610.000 4.000 610.600 ;
    END
  END vb_din0[29]
  PIN vb_din0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 87.760 4.000 88.360 ;
    END
  END vb_din0[2]
  PIN vb_din0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 624.960 4.000 625.560 ;
    END
  END vb_din0[30]
  PIN vb_din0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 640.600 4.000 641.200 ;
    END
  END vb_din0[31]
  PIN vb_din0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 118.360 4.000 118.960 ;
    END
  END vb_din0[3]
  PIN vb_din0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 148.960 4.000 149.560 ;
    END
  END vb_din0[4]
  PIN vb_din0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 174.120 4.000 174.720 ;
    END
  END vb_din0[5]
  PIN vb_din0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 199.280 4.000 199.880 ;
    END
  END vb_din0[6]
  PIN vb_din0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 224.440 4.000 225.040 ;
    END
  END vb_din0[7]
  PIN vb_din0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 250.280 4.000 250.880 ;
    END
  END vb_din0[8]
  PIN vb_din0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 275.440 4.000 276.040 ;
    END
  END vb_din0[9]
  PIN vb_dout0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.000 4.000 32.600 ;
    END
  END vb_dout0[0]
  PIN vb_dout0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 306.040 4.000 306.640 ;
    END
  END vb_dout0[10]
  PIN vb_dout0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 331.200 4.000 331.800 ;
    END
  END vb_dout0[11]
  PIN vb_dout0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 356.360 4.000 356.960 ;
    END
  END vb_dout0[12]
  PIN vb_dout0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 372.000 4.000 372.600 ;
    END
  END vb_dout0[13]
  PIN vb_dout0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 386.960 4.000 387.560 ;
    END
  END vb_dout0[14]
  PIN vb_dout0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 401.920 4.000 402.520 ;
    END
  END vb_dout0[15]
  PIN vb_dout0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 417.560 4.000 418.160 ;
    END
  END vb_dout0[16]
  PIN vb_dout0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 432.520 4.000 433.120 ;
    END
  END vb_dout0[17]
  PIN vb_dout0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 447.480 4.000 448.080 ;
    END
  END vb_dout0[18]
  PIN vb_dout0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 463.120 4.000 463.720 ;
    END
  END vb_dout0[19]
  PIN vb_dout0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 62.600 4.000 63.200 ;
    END
  END vb_dout0[1]
  PIN vb_dout0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 478.080 4.000 478.680 ;
    END
  END vb_dout0[20]
  PIN vb_dout0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 493.040 4.000 493.640 ;
    END
  END vb_dout0[21]
  PIN vb_dout0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 508.680 4.000 509.280 ;
    END
  END vb_dout0[22]
  PIN vb_dout0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 523.640 4.000 524.240 ;
    END
  END vb_dout0[23]
  PIN vb_dout0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 538.600 4.000 539.200 ;
    END
  END vb_dout0[24]
  PIN vb_dout0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 554.240 4.000 554.840 ;
    END
  END vb_dout0[25]
  PIN vb_dout0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 569.200 4.000 569.800 ;
    END
  END vb_dout0[26]
  PIN vb_dout0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 584.840 4.000 585.440 ;
    END
  END vb_dout0[27]
  PIN vb_dout0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 599.800 4.000 600.400 ;
    END
  END vb_dout0[28]
  PIN vb_dout0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 614.760 4.000 615.360 ;
    END
  END vb_dout0[29]
  PIN vb_dout0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.200 4.000 93.800 ;
    END
  END vb_dout0[2]
  PIN vb_dout0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 630.400 4.000 631.000 ;
    END
  END vb_dout0[30]
  PIN vb_dout0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 645.360 4.000 645.960 ;
    END
  END vb_dout0[31]
  PIN vb_dout0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 123.120 4.000 123.720 ;
    END
  END vb_dout0[3]
  PIN vb_dout0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.720 4.000 154.320 ;
    END
  END vb_dout0[4]
  PIN vb_dout0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 178.880 4.000 179.480 ;
    END
  END vb_dout0[5]
  PIN vb_dout0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.720 4.000 205.320 ;
    END
  END vb_dout0[6]
  PIN vb_dout0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 229.880 4.000 230.480 ;
    END
  END vb_dout0[7]
  PIN vb_dout0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 255.040 4.000 255.640 ;
    END
  END vb_dout0[8]
  PIN vb_dout0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 280.200 4.000 280.800 ;
    END
  END vb_dout0[9]
  PIN vb_dout1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END vb_dout1[0]
  PIN vb_dout1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 310.800 4.000 311.400 ;
    END
  END vb_dout1[10]
  PIN vb_dout1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 335.960 4.000 336.560 ;
    END
  END vb_dout1[11]
  PIN vb_dout1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 361.800 4.000 362.400 ;
    END
  END vb_dout1[12]
  PIN vb_dout1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 376.760 4.000 377.360 ;
    END
  END vb_dout1[13]
  PIN vb_dout1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 391.720 4.000 392.320 ;
    END
  END vb_dout1[14]
  PIN vb_dout1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 407.360 4.000 407.960 ;
    END
  END vb_dout1[15]
  PIN vb_dout1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 422.320 4.000 422.920 ;
    END
  END vb_dout1[16]
  PIN vb_dout1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 437.280 4.000 437.880 ;
    END
  END vb_dout1[17]
  PIN vb_dout1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 452.920 4.000 453.520 ;
    END
  END vb_dout1[18]
  PIN vb_dout1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 467.880 4.000 468.480 ;
    END
  END vb_dout1[19]
  PIN vb_dout1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 67.360 4.000 67.960 ;
    END
  END vb_dout1[1]
  PIN vb_dout1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 483.520 4.000 484.120 ;
    END
  END vb_dout1[20]
  PIN vb_dout1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 498.480 4.000 499.080 ;
    END
  END vb_dout1[21]
  PIN vb_dout1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 513.440 4.000 514.040 ;
    END
  END vb_dout1[22]
  PIN vb_dout1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 529.080 4.000 529.680 ;
    END
  END vb_dout1[23]
  PIN vb_dout1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 544.040 4.000 544.640 ;
    END
  END vb_dout1[24]
  PIN vb_dout1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 559.000 4.000 559.600 ;
    END
  END vb_dout1[25]
  PIN vb_dout1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 574.640 4.000 575.240 ;
    END
  END vb_dout1[26]
  PIN vb_dout1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 589.600 4.000 590.200 ;
    END
  END vb_dout1[27]
  PIN vb_dout1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 604.560 4.000 605.160 ;
    END
  END vb_dout1[28]
  PIN vb_dout1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 620.200 4.000 620.800 ;
    END
  END vb_dout1[29]
  PIN vb_dout1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 97.960 4.000 98.560 ;
    END
  END vb_dout1[2]
  PIN vb_dout1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 635.160 4.000 635.760 ;
    END
  END vb_dout1[30]
  PIN vb_dout1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 650.120 4.000 650.720 ;
    END
  END vb_dout1[31]
  PIN vb_dout1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 128.560 4.000 129.160 ;
    END
  END vb_dout1[3]
  PIN vb_dout1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.160 4.000 159.760 ;
    END
  END vb_dout1[4]
  PIN vb_dout1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 184.320 4.000 184.920 ;
    END
  END vb_dout1[5]
  PIN vb_dout1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 209.480 4.000 210.080 ;
    END
  END vb_dout1[6]
  PIN vb_dout1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 234.640 4.000 235.240 ;
    END
  END vb_dout1[7]
  PIN vb_dout1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 260.480 4.000 261.080 ;
    END
  END vb_dout1[8]
  PIN vb_dout1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 285.640 4.000 286.240 ;
    END
  END vb_dout1[9]
  PIN vb_web0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 11.600 4.000 12.200 ;
    END
  END vb_web0
  PIN vb_wmask0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.200 4.000 42.800 ;
    END
  END vb_wmask0[0]
  PIN vb_wmask0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.800 4.000 73.400 ;
    END
  END vb_wmask0[1]
  PIN vb_wmask0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 103.400 4.000 104.000 ;
    END
  END vb_wmask0[2]
  PIN vb_wmask0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 133.320 4.000 133.920 ;
    END
  END vb_wmask0[3]
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.840 10.640 1251.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1403.440 10.640 1405.040 1488.080 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1326.640 10.640 1328.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1480.240 10.640 1481.840 1488.080 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 1494.080 1487.925 ;
      LAYER met1 ;
        RECT 2.370 9.900 1494.080 1488.080 ;
      LAYER met2 ;
        RECT 2.400 4.280 1489.840 1497.205 ;
        RECT 2.400 2.195 9.470 4.280 ;
        RECT 10.310 2.195 29.250 4.280 ;
        RECT 30.090 2.195 49.030 4.280 ;
        RECT 49.870 2.195 69.270 4.280 ;
        RECT 70.110 2.195 89.050 4.280 ;
        RECT 89.890 2.195 109.290 4.280 ;
        RECT 110.130 2.195 129.070 4.280 ;
        RECT 129.910 2.195 149.310 4.280 ;
        RECT 150.150 2.195 169.090 4.280 ;
        RECT 169.930 2.195 189.330 4.280 ;
        RECT 190.170 2.195 209.110 4.280 ;
        RECT 209.950 2.195 229.350 4.280 ;
        RECT 230.190 2.195 249.130 4.280 ;
        RECT 249.970 2.195 269.370 4.280 ;
        RECT 270.210 2.195 289.150 4.280 ;
        RECT 289.990 2.195 309.390 4.280 ;
        RECT 310.230 2.195 329.170 4.280 ;
        RECT 330.010 2.195 349.410 4.280 ;
        RECT 350.250 2.195 369.190 4.280 ;
        RECT 370.030 2.195 389.430 4.280 ;
        RECT 390.270 2.195 409.210 4.280 ;
        RECT 410.050 2.195 429.450 4.280 ;
        RECT 430.290 2.195 449.230 4.280 ;
        RECT 450.070 2.195 469.470 4.280 ;
        RECT 470.310 2.195 489.250 4.280 ;
        RECT 490.090 2.195 509.490 4.280 ;
        RECT 510.330 2.195 529.270 4.280 ;
        RECT 530.110 2.195 549.050 4.280 ;
        RECT 549.890 2.195 569.290 4.280 ;
        RECT 570.130 2.195 589.070 4.280 ;
        RECT 589.910 2.195 609.310 4.280 ;
        RECT 610.150 2.195 629.090 4.280 ;
        RECT 629.930 2.195 649.330 4.280 ;
        RECT 650.170 2.195 669.110 4.280 ;
        RECT 669.950 2.195 689.350 4.280 ;
        RECT 690.190 2.195 709.130 4.280 ;
        RECT 709.970 2.195 729.370 4.280 ;
        RECT 730.210 2.195 749.150 4.280 ;
        RECT 749.990 2.195 769.390 4.280 ;
        RECT 770.230 2.195 789.170 4.280 ;
        RECT 790.010 2.195 809.410 4.280 ;
        RECT 810.250 2.195 829.190 4.280 ;
        RECT 830.030 2.195 849.430 4.280 ;
        RECT 850.270 2.195 869.210 4.280 ;
        RECT 870.050 2.195 889.450 4.280 ;
        RECT 890.290 2.195 909.230 4.280 ;
        RECT 910.070 2.195 929.470 4.280 ;
        RECT 930.310 2.195 949.250 4.280 ;
        RECT 950.090 2.195 969.490 4.280 ;
        RECT 970.330 2.195 989.270 4.280 ;
        RECT 990.110 2.195 1009.510 4.280 ;
        RECT 1010.350 2.195 1029.290 4.280 ;
        RECT 1030.130 2.195 1049.070 4.280 ;
        RECT 1049.910 2.195 1069.310 4.280 ;
        RECT 1070.150 2.195 1089.090 4.280 ;
        RECT 1089.930 2.195 1109.330 4.280 ;
        RECT 1110.170 2.195 1129.110 4.280 ;
        RECT 1129.950 2.195 1149.350 4.280 ;
        RECT 1150.190 2.195 1169.130 4.280 ;
        RECT 1169.970 2.195 1189.370 4.280 ;
        RECT 1190.210 2.195 1209.150 4.280 ;
        RECT 1209.990 2.195 1229.390 4.280 ;
        RECT 1230.230 2.195 1249.170 4.280 ;
        RECT 1250.010 2.195 1269.410 4.280 ;
        RECT 1270.250 2.195 1289.190 4.280 ;
        RECT 1290.030 2.195 1309.430 4.280 ;
        RECT 1310.270 2.195 1329.210 4.280 ;
        RECT 1330.050 2.195 1349.450 4.280 ;
        RECT 1350.290 2.195 1369.230 4.280 ;
        RECT 1370.070 2.195 1389.470 4.280 ;
        RECT 1390.310 2.195 1409.250 4.280 ;
        RECT 1410.090 2.195 1429.490 4.280 ;
        RECT 1430.330 2.195 1449.270 4.280 ;
        RECT 1450.110 2.195 1469.510 4.280 ;
        RECT 1470.350 2.195 1489.290 4.280 ;
      LAYER met3 ;
        RECT 4.400 1496.320 1481.840 1497.185 ;
        RECT 4.000 1492.960 1481.840 1496.320 ;
        RECT 4.400 1491.560 1481.840 1492.960 ;
        RECT 4.000 1487.520 1481.840 1491.560 ;
        RECT 4.400 1486.120 1481.840 1487.520 ;
        RECT 4.000 1482.760 1481.840 1486.120 ;
        RECT 4.400 1481.360 1481.840 1482.760 ;
        RECT 4.000 1477.320 1481.840 1481.360 ;
        RECT 4.400 1475.920 1481.840 1477.320 ;
        RECT 4.000 1472.560 1481.840 1475.920 ;
        RECT 4.400 1471.160 1481.840 1472.560 ;
        RECT 4.000 1467.120 1481.840 1471.160 ;
        RECT 4.400 1465.720 1481.840 1467.120 ;
        RECT 4.000 1462.360 1481.840 1465.720 ;
        RECT 4.400 1460.960 1481.840 1462.360 ;
        RECT 4.000 1456.920 1481.840 1460.960 ;
        RECT 4.400 1455.520 1481.840 1456.920 ;
        RECT 4.000 1452.160 1481.840 1455.520 ;
        RECT 4.400 1450.760 1481.840 1452.160 ;
        RECT 4.000 1447.400 1481.840 1450.760 ;
        RECT 4.400 1446.000 1481.840 1447.400 ;
        RECT 4.000 1441.960 1481.840 1446.000 ;
        RECT 4.400 1440.560 1481.840 1441.960 ;
        RECT 4.000 1437.200 1481.840 1440.560 ;
        RECT 4.400 1435.800 1481.840 1437.200 ;
        RECT 4.000 1431.760 1481.840 1435.800 ;
        RECT 4.400 1430.360 1481.840 1431.760 ;
        RECT 4.000 1427.000 1481.840 1430.360 ;
        RECT 4.400 1425.600 1481.840 1427.000 ;
        RECT 4.000 1421.560 1481.840 1425.600 ;
        RECT 4.400 1420.160 1481.840 1421.560 ;
        RECT 4.000 1416.800 1481.840 1420.160 ;
        RECT 4.400 1415.400 1481.840 1416.800 ;
        RECT 4.000 1411.360 1481.840 1415.400 ;
        RECT 4.400 1409.960 1481.840 1411.360 ;
        RECT 4.000 1406.600 1481.840 1409.960 ;
        RECT 4.400 1405.200 1481.840 1406.600 ;
        RECT 4.000 1401.160 1481.840 1405.200 ;
        RECT 4.400 1399.760 1481.840 1401.160 ;
        RECT 4.000 1396.400 1481.840 1399.760 ;
        RECT 4.400 1395.000 1481.840 1396.400 ;
        RECT 4.000 1391.640 1481.840 1395.000 ;
        RECT 4.400 1390.240 1481.840 1391.640 ;
        RECT 4.000 1386.200 1481.840 1390.240 ;
        RECT 4.400 1384.800 1481.840 1386.200 ;
        RECT 4.000 1381.440 1481.840 1384.800 ;
        RECT 4.400 1380.040 1481.840 1381.440 ;
        RECT 4.000 1376.000 1481.840 1380.040 ;
        RECT 4.400 1374.600 1481.840 1376.000 ;
        RECT 4.000 1371.240 1481.840 1374.600 ;
        RECT 4.400 1369.840 1481.840 1371.240 ;
        RECT 4.000 1365.800 1481.840 1369.840 ;
        RECT 4.400 1364.400 1481.840 1365.800 ;
        RECT 4.000 1361.040 1481.840 1364.400 ;
        RECT 4.400 1359.640 1481.840 1361.040 ;
        RECT 4.000 1355.600 1481.840 1359.640 ;
        RECT 4.400 1354.200 1481.840 1355.600 ;
        RECT 4.000 1350.840 1481.840 1354.200 ;
        RECT 4.400 1349.440 1481.840 1350.840 ;
        RECT 4.000 1345.400 1481.840 1349.440 ;
        RECT 4.400 1344.000 1481.840 1345.400 ;
        RECT 4.000 1340.640 1481.840 1344.000 ;
        RECT 4.400 1339.240 1481.840 1340.640 ;
        RECT 4.000 1335.880 1481.840 1339.240 ;
        RECT 4.400 1334.480 1481.840 1335.880 ;
        RECT 4.000 1330.440 1481.840 1334.480 ;
        RECT 4.400 1329.040 1481.840 1330.440 ;
        RECT 4.000 1325.680 1481.840 1329.040 ;
        RECT 4.400 1324.280 1481.840 1325.680 ;
        RECT 4.000 1320.240 1481.840 1324.280 ;
        RECT 4.400 1318.840 1481.840 1320.240 ;
        RECT 4.000 1315.480 1481.840 1318.840 ;
        RECT 4.400 1314.080 1481.840 1315.480 ;
        RECT 4.000 1310.040 1481.840 1314.080 ;
        RECT 4.400 1308.640 1481.840 1310.040 ;
        RECT 4.000 1305.280 1481.840 1308.640 ;
        RECT 4.400 1303.880 1481.840 1305.280 ;
        RECT 4.000 1299.840 1481.840 1303.880 ;
        RECT 4.400 1298.440 1481.840 1299.840 ;
        RECT 4.000 1295.080 1481.840 1298.440 ;
        RECT 4.400 1293.680 1481.840 1295.080 ;
        RECT 4.000 1289.640 1481.840 1293.680 ;
        RECT 4.400 1288.240 1481.840 1289.640 ;
        RECT 4.000 1284.880 1481.840 1288.240 ;
        RECT 4.400 1283.480 1481.840 1284.880 ;
        RECT 4.000 1280.120 1481.840 1283.480 ;
        RECT 4.400 1278.720 1481.840 1280.120 ;
        RECT 4.000 1274.680 1481.840 1278.720 ;
        RECT 4.400 1273.280 1481.840 1274.680 ;
        RECT 4.000 1269.920 1481.840 1273.280 ;
        RECT 4.400 1268.520 1481.840 1269.920 ;
        RECT 4.000 1264.480 1481.840 1268.520 ;
        RECT 4.400 1263.080 1481.840 1264.480 ;
        RECT 4.000 1259.720 1481.840 1263.080 ;
        RECT 4.400 1258.320 1481.840 1259.720 ;
        RECT 4.000 1254.280 1481.840 1258.320 ;
        RECT 4.400 1252.880 1481.840 1254.280 ;
        RECT 4.000 1249.520 1481.840 1252.880 ;
        RECT 4.400 1248.120 1481.840 1249.520 ;
        RECT 4.000 1244.080 1481.840 1248.120 ;
        RECT 4.400 1242.680 1481.840 1244.080 ;
        RECT 4.000 1239.320 1481.840 1242.680 ;
        RECT 4.400 1237.920 1481.840 1239.320 ;
        RECT 4.000 1234.560 1481.840 1237.920 ;
        RECT 4.400 1233.160 1481.840 1234.560 ;
        RECT 4.000 1229.120 1481.840 1233.160 ;
        RECT 4.400 1227.720 1481.840 1229.120 ;
        RECT 4.000 1224.360 1481.840 1227.720 ;
        RECT 4.400 1222.960 1481.840 1224.360 ;
        RECT 4.000 1218.920 1481.840 1222.960 ;
        RECT 4.400 1217.520 1481.840 1218.920 ;
        RECT 4.000 1214.160 1481.840 1217.520 ;
        RECT 4.400 1212.760 1481.840 1214.160 ;
        RECT 4.000 1208.720 1481.840 1212.760 ;
        RECT 4.400 1207.320 1481.840 1208.720 ;
        RECT 4.000 1203.960 1481.840 1207.320 ;
        RECT 4.400 1202.560 1481.840 1203.960 ;
        RECT 4.000 1198.520 1481.840 1202.560 ;
        RECT 4.400 1197.120 1481.840 1198.520 ;
        RECT 4.000 1193.760 1481.840 1197.120 ;
        RECT 4.400 1192.360 1481.840 1193.760 ;
        RECT 4.000 1188.320 1481.840 1192.360 ;
        RECT 4.400 1186.920 1481.840 1188.320 ;
        RECT 4.000 1183.560 1481.840 1186.920 ;
        RECT 4.400 1182.160 1481.840 1183.560 ;
        RECT 4.000 1178.800 1481.840 1182.160 ;
        RECT 4.400 1177.400 1481.840 1178.800 ;
        RECT 4.000 1173.360 1481.840 1177.400 ;
        RECT 4.400 1171.960 1481.840 1173.360 ;
        RECT 4.000 1168.600 1481.840 1171.960 ;
        RECT 4.400 1167.200 1481.840 1168.600 ;
        RECT 4.000 1163.160 1481.840 1167.200 ;
        RECT 4.400 1161.760 1481.840 1163.160 ;
        RECT 4.000 1158.400 1481.840 1161.760 ;
        RECT 4.400 1157.000 1481.840 1158.400 ;
        RECT 4.000 1152.960 1481.840 1157.000 ;
        RECT 4.400 1151.560 1481.840 1152.960 ;
        RECT 4.000 1148.200 1481.840 1151.560 ;
        RECT 4.400 1146.800 1481.840 1148.200 ;
        RECT 4.000 1142.760 1481.840 1146.800 ;
        RECT 4.400 1141.360 1481.840 1142.760 ;
        RECT 4.000 1138.000 1481.840 1141.360 ;
        RECT 4.400 1136.600 1481.840 1138.000 ;
        RECT 4.000 1132.560 1481.840 1136.600 ;
        RECT 4.400 1131.160 1481.840 1132.560 ;
        RECT 4.000 1127.800 1481.840 1131.160 ;
        RECT 4.400 1126.400 1481.840 1127.800 ;
        RECT 4.000 1123.040 1481.840 1126.400 ;
        RECT 4.400 1121.640 1481.840 1123.040 ;
        RECT 4.000 1117.600 1481.840 1121.640 ;
        RECT 4.400 1116.200 1481.840 1117.600 ;
        RECT 4.000 1112.840 1481.840 1116.200 ;
        RECT 4.400 1111.440 1481.840 1112.840 ;
        RECT 4.000 1107.400 1481.840 1111.440 ;
        RECT 4.400 1106.000 1481.840 1107.400 ;
        RECT 4.000 1102.640 1481.840 1106.000 ;
        RECT 4.400 1101.240 1481.840 1102.640 ;
        RECT 4.000 1097.200 1481.840 1101.240 ;
        RECT 4.400 1095.800 1481.840 1097.200 ;
        RECT 4.000 1092.440 1481.840 1095.800 ;
        RECT 4.400 1091.040 1481.840 1092.440 ;
        RECT 4.000 1087.000 1481.840 1091.040 ;
        RECT 4.400 1085.600 1481.840 1087.000 ;
        RECT 4.000 1082.240 1481.840 1085.600 ;
        RECT 4.400 1080.840 1481.840 1082.240 ;
        RECT 4.000 1076.800 1481.840 1080.840 ;
        RECT 4.400 1075.400 1481.840 1076.800 ;
        RECT 4.000 1072.040 1481.840 1075.400 ;
        RECT 4.400 1070.640 1481.840 1072.040 ;
        RECT 4.000 1067.280 1481.840 1070.640 ;
        RECT 4.400 1065.880 1481.840 1067.280 ;
        RECT 4.000 1061.840 1481.840 1065.880 ;
        RECT 4.400 1060.440 1481.840 1061.840 ;
        RECT 4.000 1057.080 1481.840 1060.440 ;
        RECT 4.400 1055.680 1481.840 1057.080 ;
        RECT 4.000 1051.640 1481.840 1055.680 ;
        RECT 4.400 1050.240 1481.840 1051.640 ;
        RECT 4.000 1046.880 1481.840 1050.240 ;
        RECT 4.400 1045.480 1481.840 1046.880 ;
        RECT 4.000 1041.440 1481.840 1045.480 ;
        RECT 4.400 1040.040 1481.840 1041.440 ;
        RECT 4.000 1036.680 1481.840 1040.040 ;
        RECT 4.400 1035.280 1481.840 1036.680 ;
        RECT 4.000 1031.240 1481.840 1035.280 ;
        RECT 4.400 1029.840 1481.840 1031.240 ;
        RECT 4.000 1026.480 1481.840 1029.840 ;
        RECT 4.400 1025.080 1481.840 1026.480 ;
        RECT 4.000 1021.040 1481.840 1025.080 ;
        RECT 4.400 1019.640 1481.840 1021.040 ;
        RECT 4.000 1016.280 1481.840 1019.640 ;
        RECT 4.400 1014.880 1481.840 1016.280 ;
        RECT 4.000 1011.520 1481.840 1014.880 ;
        RECT 4.400 1010.120 1481.840 1011.520 ;
        RECT 4.000 1006.080 1481.840 1010.120 ;
        RECT 4.400 1004.680 1481.840 1006.080 ;
        RECT 4.000 1001.320 1481.840 1004.680 ;
        RECT 4.400 999.920 1481.840 1001.320 ;
        RECT 4.000 995.880 1481.840 999.920 ;
        RECT 4.400 994.480 1481.840 995.880 ;
        RECT 4.000 991.120 1481.840 994.480 ;
        RECT 4.400 989.720 1481.840 991.120 ;
        RECT 4.000 985.680 1481.840 989.720 ;
        RECT 4.400 984.280 1481.840 985.680 ;
        RECT 4.000 980.920 1481.840 984.280 ;
        RECT 4.400 979.520 1481.840 980.920 ;
        RECT 4.000 975.480 1481.840 979.520 ;
        RECT 4.400 974.080 1481.840 975.480 ;
        RECT 4.000 970.720 1481.840 974.080 ;
        RECT 4.400 969.320 1481.840 970.720 ;
        RECT 4.000 965.960 1481.840 969.320 ;
        RECT 4.400 964.560 1481.840 965.960 ;
        RECT 4.000 960.520 1481.840 964.560 ;
        RECT 4.400 959.120 1481.840 960.520 ;
        RECT 4.000 955.760 1481.840 959.120 ;
        RECT 4.400 954.360 1481.840 955.760 ;
        RECT 4.000 950.320 1481.840 954.360 ;
        RECT 4.400 948.920 1481.840 950.320 ;
        RECT 4.000 945.560 1481.840 948.920 ;
        RECT 4.400 944.160 1481.840 945.560 ;
        RECT 4.000 940.120 1481.840 944.160 ;
        RECT 4.400 938.720 1481.840 940.120 ;
        RECT 4.000 935.360 1481.840 938.720 ;
        RECT 4.400 933.960 1481.840 935.360 ;
        RECT 4.000 929.920 1481.840 933.960 ;
        RECT 4.400 928.520 1481.840 929.920 ;
        RECT 4.000 925.160 1481.840 928.520 ;
        RECT 4.400 923.760 1481.840 925.160 ;
        RECT 4.000 919.720 1481.840 923.760 ;
        RECT 4.400 918.320 1481.840 919.720 ;
        RECT 4.000 914.960 1481.840 918.320 ;
        RECT 4.400 913.560 1481.840 914.960 ;
        RECT 4.000 910.200 1481.840 913.560 ;
        RECT 4.400 908.800 1481.840 910.200 ;
        RECT 4.000 904.760 1481.840 908.800 ;
        RECT 4.400 903.360 1481.840 904.760 ;
        RECT 4.000 900.000 1481.840 903.360 ;
        RECT 4.400 898.600 1481.840 900.000 ;
        RECT 4.000 894.560 1481.840 898.600 ;
        RECT 4.400 893.160 1481.840 894.560 ;
        RECT 4.000 889.800 1481.840 893.160 ;
        RECT 4.400 888.400 1481.840 889.800 ;
        RECT 4.000 884.360 1481.840 888.400 ;
        RECT 4.400 882.960 1481.840 884.360 ;
        RECT 4.000 879.600 1481.840 882.960 ;
        RECT 4.400 878.200 1481.840 879.600 ;
        RECT 4.000 874.160 1481.840 878.200 ;
        RECT 4.400 872.760 1481.840 874.160 ;
        RECT 4.000 869.400 1481.840 872.760 ;
        RECT 4.400 868.000 1481.840 869.400 ;
        RECT 4.000 863.960 1481.840 868.000 ;
        RECT 4.400 862.560 1481.840 863.960 ;
        RECT 4.000 859.200 1481.840 862.560 ;
        RECT 4.400 857.800 1481.840 859.200 ;
        RECT 4.000 854.440 1481.840 857.800 ;
        RECT 4.400 853.040 1481.840 854.440 ;
        RECT 4.000 849.000 1481.840 853.040 ;
        RECT 4.400 847.600 1481.840 849.000 ;
        RECT 4.000 844.240 1481.840 847.600 ;
        RECT 4.400 842.840 1481.840 844.240 ;
        RECT 4.000 838.800 1481.840 842.840 ;
        RECT 4.400 837.400 1481.840 838.800 ;
        RECT 4.000 834.040 1481.840 837.400 ;
        RECT 4.400 832.640 1481.840 834.040 ;
        RECT 4.000 828.600 1481.840 832.640 ;
        RECT 4.400 827.200 1481.840 828.600 ;
        RECT 4.000 823.840 1481.840 827.200 ;
        RECT 4.400 822.440 1481.840 823.840 ;
        RECT 4.000 818.400 1481.840 822.440 ;
        RECT 4.400 817.000 1481.840 818.400 ;
        RECT 4.000 813.640 1481.840 817.000 ;
        RECT 4.400 812.240 1481.840 813.640 ;
        RECT 4.000 808.200 1481.840 812.240 ;
        RECT 4.400 806.800 1481.840 808.200 ;
        RECT 4.000 803.440 1481.840 806.800 ;
        RECT 4.400 802.040 1481.840 803.440 ;
        RECT 4.000 798.680 1481.840 802.040 ;
        RECT 4.400 797.280 1481.840 798.680 ;
        RECT 4.000 793.240 1481.840 797.280 ;
        RECT 4.400 791.840 1481.840 793.240 ;
        RECT 4.000 788.480 1481.840 791.840 ;
        RECT 4.400 787.080 1481.840 788.480 ;
        RECT 4.000 783.040 1481.840 787.080 ;
        RECT 4.400 781.640 1481.840 783.040 ;
        RECT 4.000 778.280 1481.840 781.640 ;
        RECT 4.400 776.880 1481.840 778.280 ;
        RECT 4.000 772.840 1481.840 776.880 ;
        RECT 4.400 771.440 1481.840 772.840 ;
        RECT 4.000 768.080 1481.840 771.440 ;
        RECT 4.400 766.680 1481.840 768.080 ;
        RECT 4.000 762.640 1481.840 766.680 ;
        RECT 4.400 761.240 1481.840 762.640 ;
        RECT 4.000 757.880 1481.840 761.240 ;
        RECT 4.400 756.480 1481.840 757.880 ;
        RECT 4.000 753.120 1481.840 756.480 ;
        RECT 4.400 751.720 1481.840 753.120 ;
        RECT 4.000 747.680 1481.840 751.720 ;
        RECT 4.400 746.280 1481.840 747.680 ;
        RECT 4.000 742.920 1481.840 746.280 ;
        RECT 4.400 741.520 1481.840 742.920 ;
        RECT 4.000 737.480 1481.840 741.520 ;
        RECT 4.400 736.080 1481.840 737.480 ;
        RECT 4.000 732.720 1481.840 736.080 ;
        RECT 4.400 731.320 1481.840 732.720 ;
        RECT 4.000 727.280 1481.840 731.320 ;
        RECT 4.400 725.880 1481.840 727.280 ;
        RECT 4.000 722.520 1481.840 725.880 ;
        RECT 4.400 721.120 1481.840 722.520 ;
        RECT 4.000 717.080 1481.840 721.120 ;
        RECT 4.400 715.680 1481.840 717.080 ;
        RECT 4.000 712.320 1481.840 715.680 ;
        RECT 4.400 710.920 1481.840 712.320 ;
        RECT 4.000 706.880 1481.840 710.920 ;
        RECT 4.400 705.480 1481.840 706.880 ;
        RECT 4.000 702.120 1481.840 705.480 ;
        RECT 4.400 700.720 1481.840 702.120 ;
        RECT 4.000 697.360 1481.840 700.720 ;
        RECT 4.400 695.960 1481.840 697.360 ;
        RECT 4.000 691.920 1481.840 695.960 ;
        RECT 4.400 690.520 1481.840 691.920 ;
        RECT 4.000 687.160 1481.840 690.520 ;
        RECT 4.400 685.760 1481.840 687.160 ;
        RECT 4.000 681.720 1481.840 685.760 ;
        RECT 4.400 680.320 1481.840 681.720 ;
        RECT 4.000 676.960 1481.840 680.320 ;
        RECT 4.400 675.560 1481.840 676.960 ;
        RECT 4.000 671.520 1481.840 675.560 ;
        RECT 4.400 670.120 1481.840 671.520 ;
        RECT 4.000 666.760 1481.840 670.120 ;
        RECT 4.400 665.360 1481.840 666.760 ;
        RECT 4.000 661.320 1481.840 665.360 ;
        RECT 4.400 659.920 1481.840 661.320 ;
        RECT 4.000 656.560 1481.840 659.920 ;
        RECT 4.400 655.160 1481.840 656.560 ;
        RECT 4.000 651.120 1481.840 655.160 ;
        RECT 4.400 649.720 1481.840 651.120 ;
        RECT 4.000 646.360 1481.840 649.720 ;
        RECT 4.400 644.960 1481.840 646.360 ;
        RECT 4.000 641.600 1481.840 644.960 ;
        RECT 4.400 640.200 1481.840 641.600 ;
        RECT 4.000 636.160 1481.840 640.200 ;
        RECT 4.400 634.760 1481.840 636.160 ;
        RECT 4.000 631.400 1481.840 634.760 ;
        RECT 4.400 630.000 1481.840 631.400 ;
        RECT 4.000 625.960 1481.840 630.000 ;
        RECT 4.400 624.560 1481.840 625.960 ;
        RECT 4.000 621.200 1481.840 624.560 ;
        RECT 4.400 619.800 1481.840 621.200 ;
        RECT 4.000 615.760 1481.840 619.800 ;
        RECT 4.400 614.360 1481.840 615.760 ;
        RECT 4.000 611.000 1481.840 614.360 ;
        RECT 4.400 609.600 1481.840 611.000 ;
        RECT 4.000 605.560 1481.840 609.600 ;
        RECT 4.400 604.160 1481.840 605.560 ;
        RECT 4.000 600.800 1481.840 604.160 ;
        RECT 4.400 599.400 1481.840 600.800 ;
        RECT 4.000 595.360 1481.840 599.400 ;
        RECT 4.400 593.960 1481.840 595.360 ;
        RECT 4.000 590.600 1481.840 593.960 ;
        RECT 4.400 589.200 1481.840 590.600 ;
        RECT 4.000 585.840 1481.840 589.200 ;
        RECT 4.400 584.440 1481.840 585.840 ;
        RECT 4.000 580.400 1481.840 584.440 ;
        RECT 4.400 579.000 1481.840 580.400 ;
        RECT 4.000 575.640 1481.840 579.000 ;
        RECT 4.400 574.240 1481.840 575.640 ;
        RECT 4.000 570.200 1481.840 574.240 ;
        RECT 4.400 568.800 1481.840 570.200 ;
        RECT 4.000 565.440 1481.840 568.800 ;
        RECT 4.400 564.040 1481.840 565.440 ;
        RECT 4.000 560.000 1481.840 564.040 ;
        RECT 4.400 558.600 1481.840 560.000 ;
        RECT 4.000 555.240 1481.840 558.600 ;
        RECT 4.400 553.840 1481.840 555.240 ;
        RECT 4.000 549.800 1481.840 553.840 ;
        RECT 4.400 548.400 1481.840 549.800 ;
        RECT 4.000 545.040 1481.840 548.400 ;
        RECT 4.400 543.640 1481.840 545.040 ;
        RECT 4.000 539.600 1481.840 543.640 ;
        RECT 4.400 538.200 1481.840 539.600 ;
        RECT 4.000 534.840 1481.840 538.200 ;
        RECT 4.400 533.440 1481.840 534.840 ;
        RECT 4.000 530.080 1481.840 533.440 ;
        RECT 4.400 528.680 1481.840 530.080 ;
        RECT 4.000 524.640 1481.840 528.680 ;
        RECT 4.400 523.240 1481.840 524.640 ;
        RECT 4.000 519.880 1481.840 523.240 ;
        RECT 4.400 518.480 1481.840 519.880 ;
        RECT 4.000 514.440 1481.840 518.480 ;
        RECT 4.400 513.040 1481.840 514.440 ;
        RECT 4.000 509.680 1481.840 513.040 ;
        RECT 4.400 508.280 1481.840 509.680 ;
        RECT 4.000 504.240 1481.840 508.280 ;
        RECT 4.400 502.840 1481.840 504.240 ;
        RECT 4.000 499.480 1481.840 502.840 ;
        RECT 4.400 498.080 1481.840 499.480 ;
        RECT 4.000 494.040 1481.840 498.080 ;
        RECT 4.400 492.640 1481.840 494.040 ;
        RECT 4.000 489.280 1481.840 492.640 ;
        RECT 4.400 487.880 1481.840 489.280 ;
        RECT 4.000 484.520 1481.840 487.880 ;
        RECT 4.400 483.120 1481.840 484.520 ;
        RECT 4.000 479.080 1481.840 483.120 ;
        RECT 4.400 477.680 1481.840 479.080 ;
        RECT 4.000 474.320 1481.840 477.680 ;
        RECT 4.400 472.920 1481.840 474.320 ;
        RECT 4.000 468.880 1481.840 472.920 ;
        RECT 4.400 467.480 1481.840 468.880 ;
        RECT 4.000 464.120 1481.840 467.480 ;
        RECT 4.400 462.720 1481.840 464.120 ;
        RECT 4.000 458.680 1481.840 462.720 ;
        RECT 4.400 457.280 1481.840 458.680 ;
        RECT 4.000 453.920 1481.840 457.280 ;
        RECT 4.400 452.520 1481.840 453.920 ;
        RECT 4.000 448.480 1481.840 452.520 ;
        RECT 4.400 447.080 1481.840 448.480 ;
        RECT 4.000 443.720 1481.840 447.080 ;
        RECT 4.400 442.320 1481.840 443.720 ;
        RECT 4.000 438.280 1481.840 442.320 ;
        RECT 4.400 436.880 1481.840 438.280 ;
        RECT 4.000 433.520 1481.840 436.880 ;
        RECT 4.400 432.120 1481.840 433.520 ;
        RECT 4.000 428.760 1481.840 432.120 ;
        RECT 4.400 427.360 1481.840 428.760 ;
        RECT 4.000 423.320 1481.840 427.360 ;
        RECT 4.400 421.920 1481.840 423.320 ;
        RECT 4.000 418.560 1481.840 421.920 ;
        RECT 4.400 417.160 1481.840 418.560 ;
        RECT 4.000 413.120 1481.840 417.160 ;
        RECT 4.400 411.720 1481.840 413.120 ;
        RECT 4.000 408.360 1481.840 411.720 ;
        RECT 4.400 406.960 1481.840 408.360 ;
        RECT 4.000 402.920 1481.840 406.960 ;
        RECT 4.400 401.520 1481.840 402.920 ;
        RECT 4.000 398.160 1481.840 401.520 ;
        RECT 4.400 396.760 1481.840 398.160 ;
        RECT 4.000 392.720 1481.840 396.760 ;
        RECT 4.400 391.320 1481.840 392.720 ;
        RECT 4.000 387.960 1481.840 391.320 ;
        RECT 4.400 386.560 1481.840 387.960 ;
        RECT 4.000 382.520 1481.840 386.560 ;
        RECT 4.400 381.120 1481.840 382.520 ;
        RECT 4.000 377.760 1481.840 381.120 ;
        RECT 4.400 376.360 1481.840 377.760 ;
        RECT 4.000 373.000 1481.840 376.360 ;
        RECT 4.400 371.600 1481.840 373.000 ;
        RECT 4.000 367.560 1481.840 371.600 ;
        RECT 4.400 366.160 1481.840 367.560 ;
        RECT 4.000 362.800 1481.840 366.160 ;
        RECT 4.400 361.400 1481.840 362.800 ;
        RECT 4.000 357.360 1481.840 361.400 ;
        RECT 4.400 355.960 1481.840 357.360 ;
        RECT 4.000 352.600 1481.840 355.960 ;
        RECT 4.400 351.200 1481.840 352.600 ;
        RECT 4.000 347.160 1481.840 351.200 ;
        RECT 4.400 345.760 1481.840 347.160 ;
        RECT 4.000 342.400 1481.840 345.760 ;
        RECT 4.400 341.000 1481.840 342.400 ;
        RECT 4.000 336.960 1481.840 341.000 ;
        RECT 4.400 335.560 1481.840 336.960 ;
        RECT 4.000 332.200 1481.840 335.560 ;
        RECT 4.400 330.800 1481.840 332.200 ;
        RECT 4.000 326.760 1481.840 330.800 ;
        RECT 4.400 325.360 1481.840 326.760 ;
        RECT 4.000 322.000 1481.840 325.360 ;
        RECT 4.400 320.600 1481.840 322.000 ;
        RECT 4.000 317.240 1481.840 320.600 ;
        RECT 4.400 315.840 1481.840 317.240 ;
        RECT 4.000 311.800 1481.840 315.840 ;
        RECT 4.400 310.400 1481.840 311.800 ;
        RECT 4.000 307.040 1481.840 310.400 ;
        RECT 4.400 305.640 1481.840 307.040 ;
        RECT 4.000 301.600 1481.840 305.640 ;
        RECT 4.400 300.200 1481.840 301.600 ;
        RECT 4.000 296.840 1481.840 300.200 ;
        RECT 4.400 295.440 1481.840 296.840 ;
        RECT 4.000 291.400 1481.840 295.440 ;
        RECT 4.400 290.000 1481.840 291.400 ;
        RECT 4.000 286.640 1481.840 290.000 ;
        RECT 4.400 285.240 1481.840 286.640 ;
        RECT 4.000 281.200 1481.840 285.240 ;
        RECT 4.400 279.800 1481.840 281.200 ;
        RECT 4.000 276.440 1481.840 279.800 ;
        RECT 4.400 275.040 1481.840 276.440 ;
        RECT 4.000 271.000 1481.840 275.040 ;
        RECT 4.400 269.600 1481.840 271.000 ;
        RECT 4.000 266.240 1481.840 269.600 ;
        RECT 4.400 264.840 1481.840 266.240 ;
        RECT 4.000 261.480 1481.840 264.840 ;
        RECT 4.400 260.080 1481.840 261.480 ;
        RECT 4.000 256.040 1481.840 260.080 ;
        RECT 4.400 254.640 1481.840 256.040 ;
        RECT 4.000 251.280 1481.840 254.640 ;
        RECT 4.400 249.880 1481.840 251.280 ;
        RECT 4.000 245.840 1481.840 249.880 ;
        RECT 4.400 244.440 1481.840 245.840 ;
        RECT 4.000 241.080 1481.840 244.440 ;
        RECT 4.400 239.680 1481.840 241.080 ;
        RECT 4.000 235.640 1481.840 239.680 ;
        RECT 4.400 234.240 1481.840 235.640 ;
        RECT 4.000 230.880 1481.840 234.240 ;
        RECT 4.400 229.480 1481.840 230.880 ;
        RECT 4.000 225.440 1481.840 229.480 ;
        RECT 4.400 224.040 1481.840 225.440 ;
        RECT 4.000 220.680 1481.840 224.040 ;
        RECT 4.400 219.280 1481.840 220.680 ;
        RECT 4.000 215.920 1481.840 219.280 ;
        RECT 4.400 214.520 1481.840 215.920 ;
        RECT 4.000 210.480 1481.840 214.520 ;
        RECT 4.400 209.080 1481.840 210.480 ;
        RECT 4.000 205.720 1481.840 209.080 ;
        RECT 4.400 204.320 1481.840 205.720 ;
        RECT 4.000 200.280 1481.840 204.320 ;
        RECT 4.400 198.880 1481.840 200.280 ;
        RECT 4.000 195.520 1481.840 198.880 ;
        RECT 4.400 194.120 1481.840 195.520 ;
        RECT 4.000 190.080 1481.840 194.120 ;
        RECT 4.400 188.680 1481.840 190.080 ;
        RECT 4.000 185.320 1481.840 188.680 ;
        RECT 4.400 183.920 1481.840 185.320 ;
        RECT 4.000 179.880 1481.840 183.920 ;
        RECT 4.400 178.480 1481.840 179.880 ;
        RECT 4.000 175.120 1481.840 178.480 ;
        RECT 4.400 173.720 1481.840 175.120 ;
        RECT 4.000 169.680 1481.840 173.720 ;
        RECT 4.400 168.280 1481.840 169.680 ;
        RECT 4.000 164.920 1481.840 168.280 ;
        RECT 4.400 163.520 1481.840 164.920 ;
        RECT 4.000 160.160 1481.840 163.520 ;
        RECT 4.400 158.760 1481.840 160.160 ;
        RECT 4.000 154.720 1481.840 158.760 ;
        RECT 4.400 153.320 1481.840 154.720 ;
        RECT 4.000 149.960 1481.840 153.320 ;
        RECT 4.400 148.560 1481.840 149.960 ;
        RECT 4.000 144.520 1481.840 148.560 ;
        RECT 4.400 143.120 1481.840 144.520 ;
        RECT 4.000 139.760 1481.840 143.120 ;
        RECT 4.400 138.360 1481.840 139.760 ;
        RECT 4.000 134.320 1481.840 138.360 ;
        RECT 4.400 132.920 1481.840 134.320 ;
        RECT 4.000 129.560 1481.840 132.920 ;
        RECT 4.400 128.160 1481.840 129.560 ;
        RECT 4.000 124.120 1481.840 128.160 ;
        RECT 4.400 122.720 1481.840 124.120 ;
        RECT 4.000 119.360 1481.840 122.720 ;
        RECT 4.400 117.960 1481.840 119.360 ;
        RECT 4.000 113.920 1481.840 117.960 ;
        RECT 4.400 112.520 1481.840 113.920 ;
        RECT 4.000 109.160 1481.840 112.520 ;
        RECT 4.400 107.760 1481.840 109.160 ;
        RECT 4.000 104.400 1481.840 107.760 ;
        RECT 4.400 103.000 1481.840 104.400 ;
        RECT 4.000 98.960 1481.840 103.000 ;
        RECT 4.400 97.560 1481.840 98.960 ;
        RECT 4.000 94.200 1481.840 97.560 ;
        RECT 4.400 92.800 1481.840 94.200 ;
        RECT 4.000 88.760 1481.840 92.800 ;
        RECT 4.400 87.360 1481.840 88.760 ;
        RECT 4.000 84.000 1481.840 87.360 ;
        RECT 4.400 82.600 1481.840 84.000 ;
        RECT 4.000 78.560 1481.840 82.600 ;
        RECT 4.400 77.160 1481.840 78.560 ;
        RECT 4.000 73.800 1481.840 77.160 ;
        RECT 4.400 72.400 1481.840 73.800 ;
        RECT 4.000 68.360 1481.840 72.400 ;
        RECT 4.400 66.960 1481.840 68.360 ;
        RECT 4.000 63.600 1481.840 66.960 ;
        RECT 4.400 62.200 1481.840 63.600 ;
        RECT 4.000 58.160 1481.840 62.200 ;
        RECT 4.400 56.760 1481.840 58.160 ;
        RECT 4.000 53.400 1481.840 56.760 ;
        RECT 4.400 52.000 1481.840 53.400 ;
        RECT 4.000 48.640 1481.840 52.000 ;
        RECT 4.400 47.240 1481.840 48.640 ;
        RECT 4.000 43.200 1481.840 47.240 ;
        RECT 4.400 41.800 1481.840 43.200 ;
        RECT 4.000 38.440 1481.840 41.800 ;
        RECT 4.400 37.040 1481.840 38.440 ;
        RECT 4.000 33.000 1481.840 37.040 ;
        RECT 4.400 31.600 1481.840 33.000 ;
        RECT 4.000 28.240 1481.840 31.600 ;
        RECT 4.400 26.840 1481.840 28.240 ;
        RECT 4.000 22.800 1481.840 26.840 ;
        RECT 4.400 21.400 1481.840 22.800 ;
        RECT 4.000 18.040 1481.840 21.400 ;
        RECT 4.400 16.640 1481.840 18.040 ;
        RECT 4.000 12.600 1481.840 16.640 ;
        RECT 4.400 11.200 1481.840 12.600 ;
        RECT 4.000 7.840 1481.840 11.200 ;
        RECT 4.400 6.440 1481.840 7.840 ;
        RECT 4.000 3.080 1481.840 6.440 ;
        RECT 4.400 2.215 1481.840 3.080 ;
      LAYER met4 ;
        RECT 4.895 13.095 20.640 1484.265 ;
        RECT 23.040 13.095 97.440 1484.265 ;
        RECT 99.840 13.095 174.240 1484.265 ;
        RECT 176.640 13.095 251.040 1484.265 ;
        RECT 253.440 13.095 327.840 1484.265 ;
        RECT 330.240 13.095 404.640 1484.265 ;
        RECT 407.040 13.095 481.440 1484.265 ;
        RECT 483.840 13.095 558.240 1484.265 ;
        RECT 560.640 13.095 635.040 1484.265 ;
        RECT 637.440 13.095 711.840 1484.265 ;
        RECT 714.240 13.095 788.640 1484.265 ;
        RECT 791.040 13.095 865.440 1484.265 ;
        RECT 867.840 13.095 890.265 1484.265 ;
  END
END c0_system
END LIBRARY


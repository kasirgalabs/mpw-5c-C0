magic
tech sky130A
magscale 1 2
timestamp 1647695770
<< obsli1 >>
rect 1104 2159 318872 317713
<< obsm1 >>
rect 382 1980 318872 317744
<< metal2 >>
rect 2134 0 2190 800
rect 6366 0 6422 800
rect 10598 0 10654 800
rect 14922 0 14978 800
rect 19154 0 19210 800
rect 23386 0 23442 800
rect 27710 0 27766 800
rect 31942 0 31998 800
rect 36174 0 36230 800
rect 40498 0 40554 800
rect 44730 0 44786 800
rect 49054 0 49110 800
rect 53286 0 53342 800
rect 57518 0 57574 800
rect 61842 0 61898 800
rect 66074 0 66130 800
rect 70306 0 70362 800
rect 74630 0 74686 800
rect 78862 0 78918 800
rect 83186 0 83242 800
rect 87418 0 87474 800
rect 91650 0 91706 800
rect 95974 0 96030 800
rect 100206 0 100262 800
rect 104438 0 104494 800
rect 108762 0 108818 800
rect 112994 0 113050 800
rect 117318 0 117374 800
rect 121550 0 121606 800
rect 125782 0 125838 800
rect 130106 0 130162 800
rect 134338 0 134394 800
rect 138570 0 138626 800
rect 142894 0 142950 800
rect 147126 0 147182 800
rect 151450 0 151506 800
rect 155682 0 155738 800
rect 159914 0 159970 800
rect 164238 0 164294 800
rect 168470 0 168526 800
rect 172702 0 172758 800
rect 177026 0 177082 800
rect 181258 0 181314 800
rect 185582 0 185638 800
rect 189814 0 189870 800
rect 194046 0 194102 800
rect 198370 0 198426 800
rect 202602 0 202658 800
rect 206834 0 206890 800
rect 211158 0 211214 800
rect 215390 0 215446 800
rect 219714 0 219770 800
rect 223946 0 224002 800
rect 228178 0 228234 800
rect 232502 0 232558 800
rect 236734 0 236790 800
rect 240966 0 241022 800
rect 245290 0 245346 800
rect 249522 0 249578 800
rect 253846 0 253902 800
rect 258078 0 258134 800
rect 262310 0 262366 800
rect 266634 0 266690 800
rect 270866 0 270922 800
rect 275098 0 275154 800
rect 279422 0 279478 800
rect 283654 0 283710 800
rect 287978 0 288034 800
rect 292210 0 292266 800
rect 296442 0 296498 800
rect 300766 0 300822 800
rect 304998 0 305054 800
rect 309230 0 309286 800
rect 313554 0 313610 800
rect 317786 0 317842 800
<< obsm2 >>
rect 388 856 317840 319433
rect 388 439 2078 856
rect 2246 439 6310 856
rect 6478 439 10542 856
rect 10710 439 14866 856
rect 15034 439 19098 856
rect 19266 439 23330 856
rect 23498 439 27654 856
rect 27822 439 31886 856
rect 32054 439 36118 856
rect 36286 439 40442 856
rect 40610 439 44674 856
rect 44842 439 48998 856
rect 49166 439 53230 856
rect 53398 439 57462 856
rect 57630 439 61786 856
rect 61954 439 66018 856
rect 66186 439 70250 856
rect 70418 439 74574 856
rect 74742 439 78806 856
rect 78974 439 83130 856
rect 83298 439 87362 856
rect 87530 439 91594 856
rect 91762 439 95918 856
rect 96086 439 100150 856
rect 100318 439 104382 856
rect 104550 439 108706 856
rect 108874 439 112938 856
rect 113106 439 117262 856
rect 117430 439 121494 856
rect 121662 439 125726 856
rect 125894 439 130050 856
rect 130218 439 134282 856
rect 134450 439 138514 856
rect 138682 439 142838 856
rect 143006 439 147070 856
rect 147238 439 151394 856
rect 151562 439 155626 856
rect 155794 439 159858 856
rect 160026 439 164182 856
rect 164350 439 168414 856
rect 168582 439 172646 856
rect 172814 439 176970 856
rect 177138 439 181202 856
rect 181370 439 185526 856
rect 185694 439 189758 856
rect 189926 439 193990 856
rect 194158 439 198314 856
rect 198482 439 202546 856
rect 202714 439 206778 856
rect 206946 439 211102 856
rect 211270 439 215334 856
rect 215502 439 219658 856
rect 219826 439 223890 856
rect 224058 439 228122 856
rect 228290 439 232446 856
rect 232614 439 236678 856
rect 236846 439 240910 856
rect 241078 439 245234 856
rect 245402 439 249466 856
rect 249634 439 253790 856
rect 253958 439 258022 856
rect 258190 439 262254 856
rect 262422 439 266578 856
rect 266746 439 270810 856
rect 270978 439 275042 856
rect 275210 439 279366 856
rect 279534 439 283598 856
rect 283766 439 287922 856
rect 288090 439 292154 856
rect 292322 439 296386 856
rect 296554 439 300710 856
rect 300878 439 304942 856
rect 305110 439 309174 856
rect 309342 439 313498 856
rect 313666 439 317730 856
<< metal3 >>
rect 0 319336 800 319456
rect 0 318248 800 318368
rect 0 317160 800 317280
rect 0 316072 800 316192
rect 0 314984 800 315104
rect 0 313896 800 314016
rect 0 312808 800 312928
rect 0 311720 800 311840
rect 0 310632 800 310752
rect 0 309544 800 309664
rect 0 308456 800 308576
rect 0 307368 800 307488
rect 0 306280 800 306400
rect 0 305192 800 305312
rect 0 304104 800 304224
rect 0 303016 800 303136
rect 0 301928 800 302048
rect 0 300840 800 300960
rect 0 299752 800 299872
rect 0 298800 800 298920
rect 0 297712 800 297832
rect 0 296624 800 296744
rect 0 295536 800 295656
rect 0 294448 800 294568
rect 0 293360 800 293480
rect 0 292272 800 292392
rect 0 291184 800 291304
rect 0 290096 800 290216
rect 0 289008 800 289128
rect 0 287920 800 288040
rect 0 286832 800 286952
rect 0 285744 800 285864
rect 0 284656 800 284776
rect 0 283568 800 283688
rect 0 282480 800 282600
rect 0 281392 800 281512
rect 0 280304 800 280424
rect 0 279216 800 279336
rect 0 278128 800 278248
rect 0 277176 800 277296
rect 0 276088 800 276208
rect 0 275000 800 275120
rect 0 273912 800 274032
rect 0 272824 800 272944
rect 0 271736 800 271856
rect 0 270648 800 270768
rect 0 269560 800 269680
rect 0 268472 800 268592
rect 0 267384 800 267504
rect 0 266296 800 266416
rect 0 265208 800 265328
rect 0 264120 800 264240
rect 0 263032 800 263152
rect 0 261944 800 262064
rect 0 260856 800 260976
rect 0 259768 800 259888
rect 0 258680 800 258800
rect 0 257592 800 257712
rect 0 256504 800 256624
rect 0 255552 800 255672
rect 0 254464 800 254584
rect 0 253376 800 253496
rect 0 252288 800 252408
rect 0 251200 800 251320
rect 0 250112 800 250232
rect 0 249024 800 249144
rect 0 247936 800 248056
rect 0 246848 800 246968
rect 0 245760 800 245880
rect 0 244672 800 244792
rect 0 243584 800 243704
rect 0 242496 800 242616
rect 0 241408 800 241528
rect 0 240320 800 240440
rect 0 239232 800 239352
rect 0 238144 800 238264
rect 0 237056 800 237176
rect 0 235968 800 236088
rect 0 235016 800 235136
rect 0 233928 800 234048
rect 0 232840 800 232960
rect 0 231752 800 231872
rect 0 230664 800 230784
rect 0 229576 800 229696
rect 0 228488 800 228608
rect 0 227400 800 227520
rect 0 226312 800 226432
rect 0 225224 800 225344
rect 0 224136 800 224256
rect 0 223048 800 223168
rect 0 221960 800 222080
rect 0 220872 800 220992
rect 0 219784 800 219904
rect 0 218696 800 218816
rect 0 217608 800 217728
rect 0 216520 800 216640
rect 0 215432 800 215552
rect 0 214344 800 214464
rect 0 213392 800 213512
rect 0 212304 800 212424
rect 0 211216 800 211336
rect 0 210128 800 210248
rect 0 209040 800 209160
rect 0 207952 800 208072
rect 0 206864 800 206984
rect 0 205776 800 205896
rect 0 204688 800 204808
rect 0 203600 800 203720
rect 0 202512 800 202632
rect 0 201424 800 201544
rect 0 200336 800 200456
rect 0 199248 800 199368
rect 0 198160 800 198280
rect 0 197072 800 197192
rect 0 195984 800 196104
rect 0 194896 800 195016
rect 0 193808 800 193928
rect 0 192720 800 192840
rect 0 191768 800 191888
rect 0 190680 800 190800
rect 0 189592 800 189712
rect 0 188504 800 188624
rect 0 187416 800 187536
rect 0 186328 800 186448
rect 0 185240 800 185360
rect 0 184152 800 184272
rect 0 183064 800 183184
rect 0 181976 800 182096
rect 0 180888 800 181008
rect 0 179800 800 179920
rect 0 178712 800 178832
rect 0 177624 800 177744
rect 0 176536 800 176656
rect 0 175448 800 175568
rect 0 174360 800 174480
rect 0 173272 800 173392
rect 0 172184 800 172304
rect 0 171096 800 171216
rect 0 170144 800 170264
rect 0 169056 800 169176
rect 0 167968 800 168088
rect 0 166880 800 167000
rect 0 165792 800 165912
rect 0 164704 800 164824
rect 0 163616 800 163736
rect 0 162528 800 162648
rect 0 161440 800 161560
rect 0 160352 800 160472
rect 0 159264 800 159384
rect 0 158176 800 158296
rect 0 157088 800 157208
rect 0 156000 800 156120
rect 0 154912 800 155032
rect 0 153824 800 153944
rect 0 152736 800 152856
rect 0 151648 800 151768
rect 0 150560 800 150680
rect 0 149608 800 149728
rect 0 148520 800 148640
rect 0 147432 800 147552
rect 0 146344 800 146464
rect 0 145256 800 145376
rect 0 144168 800 144288
rect 0 143080 800 143200
rect 0 141992 800 142112
rect 0 140904 800 141024
rect 0 139816 800 139936
rect 0 138728 800 138848
rect 0 137640 800 137760
rect 0 136552 800 136672
rect 0 135464 800 135584
rect 0 134376 800 134496
rect 0 133288 800 133408
rect 0 132200 800 132320
rect 0 131112 800 131232
rect 0 130024 800 130144
rect 0 128936 800 129056
rect 0 127984 800 128104
rect 0 126896 800 127016
rect 0 125808 800 125928
rect 0 124720 800 124840
rect 0 123632 800 123752
rect 0 122544 800 122664
rect 0 121456 800 121576
rect 0 120368 800 120488
rect 0 119280 800 119400
rect 0 118192 800 118312
rect 0 117104 800 117224
rect 0 116016 800 116136
rect 0 114928 800 115048
rect 0 113840 800 113960
rect 0 112752 800 112872
rect 0 111664 800 111784
rect 0 110576 800 110696
rect 0 109488 800 109608
rect 0 108400 800 108520
rect 0 107312 800 107432
rect 0 106360 800 106480
rect 0 105272 800 105392
rect 0 104184 800 104304
rect 0 103096 800 103216
rect 0 102008 800 102128
rect 0 100920 800 101040
rect 0 99832 800 99952
rect 0 98744 800 98864
rect 0 97656 800 97776
rect 0 96568 800 96688
rect 0 95480 800 95600
rect 0 94392 800 94512
rect 0 93304 800 93424
rect 0 92216 800 92336
rect 0 91128 800 91248
rect 0 90040 800 90160
rect 0 88952 800 89072
rect 0 87864 800 87984
rect 0 86776 800 86896
rect 0 85688 800 85808
rect 0 84736 800 84856
rect 0 83648 800 83768
rect 0 82560 800 82680
rect 0 81472 800 81592
rect 0 80384 800 80504
rect 0 79296 800 79416
rect 0 78208 800 78328
rect 0 77120 800 77240
rect 0 76032 800 76152
rect 0 74944 800 75064
rect 0 73856 800 73976
rect 0 72768 800 72888
rect 0 71680 800 71800
rect 0 70592 800 70712
rect 0 69504 800 69624
rect 0 68416 800 68536
rect 0 67328 800 67448
rect 0 66240 800 66360
rect 0 65152 800 65272
rect 0 64200 800 64320
rect 0 63112 800 63232
rect 0 62024 800 62144
rect 0 60936 800 61056
rect 0 59848 800 59968
rect 0 58760 800 58880
rect 0 57672 800 57792
rect 0 56584 800 56704
rect 0 55496 800 55616
rect 0 54408 800 54528
rect 0 53320 800 53440
rect 0 52232 800 52352
rect 0 51144 800 51264
rect 0 50056 800 50176
rect 0 48968 800 49088
rect 0 47880 800 48000
rect 0 46792 800 46912
rect 0 45704 800 45824
rect 0 44616 800 44736
rect 0 43528 800 43648
rect 0 42576 800 42696
rect 0 41488 800 41608
rect 0 40400 800 40520
rect 0 39312 800 39432
rect 0 38224 800 38344
rect 0 37136 800 37256
rect 0 36048 800 36168
rect 0 34960 800 35080
rect 0 33872 800 33992
rect 0 32784 800 32904
rect 0 31696 800 31816
rect 0 30608 800 30728
rect 0 29520 800 29640
rect 0 28432 800 28552
rect 0 27344 800 27464
rect 0 26256 800 26376
rect 0 25168 800 25288
rect 0 24080 800 24200
rect 0 22992 800 23112
rect 0 21904 800 22024
rect 0 20952 800 21072
rect 0 19864 800 19984
rect 0 18776 800 18896
rect 0 17688 800 17808
rect 0 16600 800 16720
rect 0 15512 800 15632
rect 0 14424 800 14544
rect 0 13336 800 13456
rect 0 12248 800 12368
rect 0 11160 800 11280
rect 0 10072 800 10192
rect 0 8984 800 9104
rect 0 7896 800 8016
rect 0 6808 800 6928
rect 0 5720 800 5840
rect 0 4632 800 4752
rect 0 3544 800 3664
rect 0 2456 800 2576
rect 0 1368 800 1488
rect 0 416 800 536
<< obsm3 >>
rect 880 319256 311728 319429
rect 800 318448 311728 319256
rect 880 318168 311728 318448
rect 800 317360 311728 318168
rect 880 317080 311728 317360
rect 800 316272 311728 317080
rect 880 315992 311728 316272
rect 800 315184 311728 315992
rect 880 314904 311728 315184
rect 800 314096 311728 314904
rect 880 313816 311728 314096
rect 800 313008 311728 313816
rect 880 312728 311728 313008
rect 800 311920 311728 312728
rect 880 311640 311728 311920
rect 800 310832 311728 311640
rect 880 310552 311728 310832
rect 800 309744 311728 310552
rect 880 309464 311728 309744
rect 800 308656 311728 309464
rect 880 308376 311728 308656
rect 800 307568 311728 308376
rect 880 307288 311728 307568
rect 800 306480 311728 307288
rect 880 306200 311728 306480
rect 800 305392 311728 306200
rect 880 305112 311728 305392
rect 800 304304 311728 305112
rect 880 304024 311728 304304
rect 800 303216 311728 304024
rect 880 302936 311728 303216
rect 800 302128 311728 302936
rect 880 301848 311728 302128
rect 800 301040 311728 301848
rect 880 300760 311728 301040
rect 800 299952 311728 300760
rect 880 299672 311728 299952
rect 800 299000 311728 299672
rect 880 298720 311728 299000
rect 800 297912 311728 298720
rect 880 297632 311728 297912
rect 800 296824 311728 297632
rect 880 296544 311728 296824
rect 800 295736 311728 296544
rect 880 295456 311728 295736
rect 800 294648 311728 295456
rect 880 294368 311728 294648
rect 800 293560 311728 294368
rect 880 293280 311728 293560
rect 800 292472 311728 293280
rect 880 292192 311728 292472
rect 800 291384 311728 292192
rect 880 291104 311728 291384
rect 800 290296 311728 291104
rect 880 290016 311728 290296
rect 800 289208 311728 290016
rect 880 288928 311728 289208
rect 800 288120 311728 288928
rect 880 287840 311728 288120
rect 800 287032 311728 287840
rect 880 286752 311728 287032
rect 800 285944 311728 286752
rect 880 285664 311728 285944
rect 800 284856 311728 285664
rect 880 284576 311728 284856
rect 800 283768 311728 284576
rect 880 283488 311728 283768
rect 800 282680 311728 283488
rect 880 282400 311728 282680
rect 800 281592 311728 282400
rect 880 281312 311728 281592
rect 800 280504 311728 281312
rect 880 280224 311728 280504
rect 800 279416 311728 280224
rect 880 279136 311728 279416
rect 800 278328 311728 279136
rect 880 278048 311728 278328
rect 800 277376 311728 278048
rect 880 277096 311728 277376
rect 800 276288 311728 277096
rect 880 276008 311728 276288
rect 800 275200 311728 276008
rect 880 274920 311728 275200
rect 800 274112 311728 274920
rect 880 273832 311728 274112
rect 800 273024 311728 273832
rect 880 272744 311728 273024
rect 800 271936 311728 272744
rect 880 271656 311728 271936
rect 800 270848 311728 271656
rect 880 270568 311728 270848
rect 800 269760 311728 270568
rect 880 269480 311728 269760
rect 800 268672 311728 269480
rect 880 268392 311728 268672
rect 800 267584 311728 268392
rect 880 267304 311728 267584
rect 800 266496 311728 267304
rect 880 266216 311728 266496
rect 800 265408 311728 266216
rect 880 265128 311728 265408
rect 800 264320 311728 265128
rect 880 264040 311728 264320
rect 800 263232 311728 264040
rect 880 262952 311728 263232
rect 800 262144 311728 262952
rect 880 261864 311728 262144
rect 800 261056 311728 261864
rect 880 260776 311728 261056
rect 800 259968 311728 260776
rect 880 259688 311728 259968
rect 800 258880 311728 259688
rect 880 258600 311728 258880
rect 800 257792 311728 258600
rect 880 257512 311728 257792
rect 800 256704 311728 257512
rect 880 256424 311728 256704
rect 800 255752 311728 256424
rect 880 255472 311728 255752
rect 800 254664 311728 255472
rect 880 254384 311728 254664
rect 800 253576 311728 254384
rect 880 253296 311728 253576
rect 800 252488 311728 253296
rect 880 252208 311728 252488
rect 800 251400 311728 252208
rect 880 251120 311728 251400
rect 800 250312 311728 251120
rect 880 250032 311728 250312
rect 800 249224 311728 250032
rect 880 248944 311728 249224
rect 800 248136 311728 248944
rect 880 247856 311728 248136
rect 800 247048 311728 247856
rect 880 246768 311728 247048
rect 800 245960 311728 246768
rect 880 245680 311728 245960
rect 800 244872 311728 245680
rect 880 244592 311728 244872
rect 800 243784 311728 244592
rect 880 243504 311728 243784
rect 800 242696 311728 243504
rect 880 242416 311728 242696
rect 800 241608 311728 242416
rect 880 241328 311728 241608
rect 800 240520 311728 241328
rect 880 240240 311728 240520
rect 800 239432 311728 240240
rect 880 239152 311728 239432
rect 800 238344 311728 239152
rect 880 238064 311728 238344
rect 800 237256 311728 238064
rect 880 236976 311728 237256
rect 800 236168 311728 236976
rect 880 235888 311728 236168
rect 800 235216 311728 235888
rect 880 234936 311728 235216
rect 800 234128 311728 234936
rect 880 233848 311728 234128
rect 800 233040 311728 233848
rect 880 232760 311728 233040
rect 800 231952 311728 232760
rect 880 231672 311728 231952
rect 800 230864 311728 231672
rect 880 230584 311728 230864
rect 800 229776 311728 230584
rect 880 229496 311728 229776
rect 800 228688 311728 229496
rect 880 228408 311728 228688
rect 800 227600 311728 228408
rect 880 227320 311728 227600
rect 800 226512 311728 227320
rect 880 226232 311728 226512
rect 800 225424 311728 226232
rect 880 225144 311728 225424
rect 800 224336 311728 225144
rect 880 224056 311728 224336
rect 800 223248 311728 224056
rect 880 222968 311728 223248
rect 800 222160 311728 222968
rect 880 221880 311728 222160
rect 800 221072 311728 221880
rect 880 220792 311728 221072
rect 800 219984 311728 220792
rect 880 219704 311728 219984
rect 800 218896 311728 219704
rect 880 218616 311728 218896
rect 800 217808 311728 218616
rect 880 217528 311728 217808
rect 800 216720 311728 217528
rect 880 216440 311728 216720
rect 800 215632 311728 216440
rect 880 215352 311728 215632
rect 800 214544 311728 215352
rect 880 214264 311728 214544
rect 800 213592 311728 214264
rect 880 213312 311728 213592
rect 800 212504 311728 213312
rect 880 212224 311728 212504
rect 800 211416 311728 212224
rect 880 211136 311728 211416
rect 800 210328 311728 211136
rect 880 210048 311728 210328
rect 800 209240 311728 210048
rect 880 208960 311728 209240
rect 800 208152 311728 208960
rect 880 207872 311728 208152
rect 800 207064 311728 207872
rect 880 206784 311728 207064
rect 800 205976 311728 206784
rect 880 205696 311728 205976
rect 800 204888 311728 205696
rect 880 204608 311728 204888
rect 800 203800 311728 204608
rect 880 203520 311728 203800
rect 800 202712 311728 203520
rect 880 202432 311728 202712
rect 800 201624 311728 202432
rect 880 201344 311728 201624
rect 800 200536 311728 201344
rect 880 200256 311728 200536
rect 800 199448 311728 200256
rect 880 199168 311728 199448
rect 800 198360 311728 199168
rect 880 198080 311728 198360
rect 800 197272 311728 198080
rect 880 196992 311728 197272
rect 800 196184 311728 196992
rect 880 195904 311728 196184
rect 800 195096 311728 195904
rect 880 194816 311728 195096
rect 800 194008 311728 194816
rect 880 193728 311728 194008
rect 800 192920 311728 193728
rect 880 192640 311728 192920
rect 800 191968 311728 192640
rect 880 191688 311728 191968
rect 800 190880 311728 191688
rect 880 190600 311728 190880
rect 800 189792 311728 190600
rect 880 189512 311728 189792
rect 800 188704 311728 189512
rect 880 188424 311728 188704
rect 800 187616 311728 188424
rect 880 187336 311728 187616
rect 800 186528 311728 187336
rect 880 186248 311728 186528
rect 800 185440 311728 186248
rect 880 185160 311728 185440
rect 800 184352 311728 185160
rect 880 184072 311728 184352
rect 800 183264 311728 184072
rect 880 182984 311728 183264
rect 800 182176 311728 182984
rect 880 181896 311728 182176
rect 800 181088 311728 181896
rect 880 180808 311728 181088
rect 800 180000 311728 180808
rect 880 179720 311728 180000
rect 800 178912 311728 179720
rect 880 178632 311728 178912
rect 800 177824 311728 178632
rect 880 177544 311728 177824
rect 800 176736 311728 177544
rect 880 176456 311728 176736
rect 800 175648 311728 176456
rect 880 175368 311728 175648
rect 800 174560 311728 175368
rect 880 174280 311728 174560
rect 800 173472 311728 174280
rect 880 173192 311728 173472
rect 800 172384 311728 173192
rect 880 172104 311728 172384
rect 800 171296 311728 172104
rect 880 171016 311728 171296
rect 800 170344 311728 171016
rect 880 170064 311728 170344
rect 800 169256 311728 170064
rect 880 168976 311728 169256
rect 800 168168 311728 168976
rect 880 167888 311728 168168
rect 800 167080 311728 167888
rect 880 166800 311728 167080
rect 800 165992 311728 166800
rect 880 165712 311728 165992
rect 800 164904 311728 165712
rect 880 164624 311728 164904
rect 800 163816 311728 164624
rect 880 163536 311728 163816
rect 800 162728 311728 163536
rect 880 162448 311728 162728
rect 800 161640 311728 162448
rect 880 161360 311728 161640
rect 800 160552 311728 161360
rect 880 160272 311728 160552
rect 800 159464 311728 160272
rect 880 159184 311728 159464
rect 800 158376 311728 159184
rect 880 158096 311728 158376
rect 800 157288 311728 158096
rect 880 157008 311728 157288
rect 800 156200 311728 157008
rect 880 155920 311728 156200
rect 800 155112 311728 155920
rect 880 154832 311728 155112
rect 800 154024 311728 154832
rect 880 153744 311728 154024
rect 800 152936 311728 153744
rect 880 152656 311728 152936
rect 800 151848 311728 152656
rect 880 151568 311728 151848
rect 800 150760 311728 151568
rect 880 150480 311728 150760
rect 800 149808 311728 150480
rect 880 149528 311728 149808
rect 800 148720 311728 149528
rect 880 148440 311728 148720
rect 800 147632 311728 148440
rect 880 147352 311728 147632
rect 800 146544 311728 147352
rect 880 146264 311728 146544
rect 800 145456 311728 146264
rect 880 145176 311728 145456
rect 800 144368 311728 145176
rect 880 144088 311728 144368
rect 800 143280 311728 144088
rect 880 143000 311728 143280
rect 800 142192 311728 143000
rect 880 141912 311728 142192
rect 800 141104 311728 141912
rect 880 140824 311728 141104
rect 800 140016 311728 140824
rect 880 139736 311728 140016
rect 800 138928 311728 139736
rect 880 138648 311728 138928
rect 800 137840 311728 138648
rect 880 137560 311728 137840
rect 800 136752 311728 137560
rect 880 136472 311728 136752
rect 800 135664 311728 136472
rect 880 135384 311728 135664
rect 800 134576 311728 135384
rect 880 134296 311728 134576
rect 800 133488 311728 134296
rect 880 133208 311728 133488
rect 800 132400 311728 133208
rect 880 132120 311728 132400
rect 800 131312 311728 132120
rect 880 131032 311728 131312
rect 800 130224 311728 131032
rect 880 129944 311728 130224
rect 800 129136 311728 129944
rect 880 128856 311728 129136
rect 800 128184 311728 128856
rect 880 127904 311728 128184
rect 800 127096 311728 127904
rect 880 126816 311728 127096
rect 800 126008 311728 126816
rect 880 125728 311728 126008
rect 800 124920 311728 125728
rect 880 124640 311728 124920
rect 800 123832 311728 124640
rect 880 123552 311728 123832
rect 800 122744 311728 123552
rect 880 122464 311728 122744
rect 800 121656 311728 122464
rect 880 121376 311728 121656
rect 800 120568 311728 121376
rect 880 120288 311728 120568
rect 800 119480 311728 120288
rect 880 119200 311728 119480
rect 800 118392 311728 119200
rect 880 118112 311728 118392
rect 800 117304 311728 118112
rect 880 117024 311728 117304
rect 800 116216 311728 117024
rect 880 115936 311728 116216
rect 800 115128 311728 115936
rect 880 114848 311728 115128
rect 800 114040 311728 114848
rect 880 113760 311728 114040
rect 800 112952 311728 113760
rect 880 112672 311728 112952
rect 800 111864 311728 112672
rect 880 111584 311728 111864
rect 800 110776 311728 111584
rect 880 110496 311728 110776
rect 800 109688 311728 110496
rect 880 109408 311728 109688
rect 800 108600 311728 109408
rect 880 108320 311728 108600
rect 800 107512 311728 108320
rect 880 107232 311728 107512
rect 800 106560 311728 107232
rect 880 106280 311728 106560
rect 800 105472 311728 106280
rect 880 105192 311728 105472
rect 800 104384 311728 105192
rect 880 104104 311728 104384
rect 800 103296 311728 104104
rect 880 103016 311728 103296
rect 800 102208 311728 103016
rect 880 101928 311728 102208
rect 800 101120 311728 101928
rect 880 100840 311728 101120
rect 800 100032 311728 100840
rect 880 99752 311728 100032
rect 800 98944 311728 99752
rect 880 98664 311728 98944
rect 800 97856 311728 98664
rect 880 97576 311728 97856
rect 800 96768 311728 97576
rect 880 96488 311728 96768
rect 800 95680 311728 96488
rect 880 95400 311728 95680
rect 800 94592 311728 95400
rect 880 94312 311728 94592
rect 800 93504 311728 94312
rect 880 93224 311728 93504
rect 800 92416 311728 93224
rect 880 92136 311728 92416
rect 800 91328 311728 92136
rect 880 91048 311728 91328
rect 800 90240 311728 91048
rect 880 89960 311728 90240
rect 800 89152 311728 89960
rect 880 88872 311728 89152
rect 800 88064 311728 88872
rect 880 87784 311728 88064
rect 800 86976 311728 87784
rect 880 86696 311728 86976
rect 800 85888 311728 86696
rect 880 85608 311728 85888
rect 800 84936 311728 85608
rect 880 84656 311728 84936
rect 800 83848 311728 84656
rect 880 83568 311728 83848
rect 800 82760 311728 83568
rect 880 82480 311728 82760
rect 800 81672 311728 82480
rect 880 81392 311728 81672
rect 800 80584 311728 81392
rect 880 80304 311728 80584
rect 800 79496 311728 80304
rect 880 79216 311728 79496
rect 800 78408 311728 79216
rect 880 78128 311728 78408
rect 800 77320 311728 78128
rect 880 77040 311728 77320
rect 800 76232 311728 77040
rect 880 75952 311728 76232
rect 800 75144 311728 75952
rect 880 74864 311728 75144
rect 800 74056 311728 74864
rect 880 73776 311728 74056
rect 800 72968 311728 73776
rect 880 72688 311728 72968
rect 800 71880 311728 72688
rect 880 71600 311728 71880
rect 800 70792 311728 71600
rect 880 70512 311728 70792
rect 800 69704 311728 70512
rect 880 69424 311728 69704
rect 800 68616 311728 69424
rect 880 68336 311728 68616
rect 800 67528 311728 68336
rect 880 67248 311728 67528
rect 800 66440 311728 67248
rect 880 66160 311728 66440
rect 800 65352 311728 66160
rect 880 65072 311728 65352
rect 800 64400 311728 65072
rect 880 64120 311728 64400
rect 800 63312 311728 64120
rect 880 63032 311728 63312
rect 800 62224 311728 63032
rect 880 61944 311728 62224
rect 800 61136 311728 61944
rect 880 60856 311728 61136
rect 800 60048 311728 60856
rect 880 59768 311728 60048
rect 800 58960 311728 59768
rect 880 58680 311728 58960
rect 800 57872 311728 58680
rect 880 57592 311728 57872
rect 800 56784 311728 57592
rect 880 56504 311728 56784
rect 800 55696 311728 56504
rect 880 55416 311728 55696
rect 800 54608 311728 55416
rect 880 54328 311728 54608
rect 800 53520 311728 54328
rect 880 53240 311728 53520
rect 800 52432 311728 53240
rect 880 52152 311728 52432
rect 800 51344 311728 52152
rect 880 51064 311728 51344
rect 800 50256 311728 51064
rect 880 49976 311728 50256
rect 800 49168 311728 49976
rect 880 48888 311728 49168
rect 800 48080 311728 48888
rect 880 47800 311728 48080
rect 800 46992 311728 47800
rect 880 46712 311728 46992
rect 800 45904 311728 46712
rect 880 45624 311728 45904
rect 800 44816 311728 45624
rect 880 44536 311728 44816
rect 800 43728 311728 44536
rect 880 43448 311728 43728
rect 800 42776 311728 43448
rect 880 42496 311728 42776
rect 800 41688 311728 42496
rect 880 41408 311728 41688
rect 800 40600 311728 41408
rect 880 40320 311728 40600
rect 800 39512 311728 40320
rect 880 39232 311728 39512
rect 800 38424 311728 39232
rect 880 38144 311728 38424
rect 800 37336 311728 38144
rect 880 37056 311728 37336
rect 800 36248 311728 37056
rect 880 35968 311728 36248
rect 800 35160 311728 35968
rect 880 34880 311728 35160
rect 800 34072 311728 34880
rect 880 33792 311728 34072
rect 800 32984 311728 33792
rect 880 32704 311728 32984
rect 800 31896 311728 32704
rect 880 31616 311728 31896
rect 800 30808 311728 31616
rect 880 30528 311728 30808
rect 800 29720 311728 30528
rect 880 29440 311728 29720
rect 800 28632 311728 29440
rect 880 28352 311728 28632
rect 800 27544 311728 28352
rect 880 27264 311728 27544
rect 800 26456 311728 27264
rect 880 26176 311728 26456
rect 800 25368 311728 26176
rect 880 25088 311728 25368
rect 800 24280 311728 25088
rect 880 24000 311728 24280
rect 800 23192 311728 24000
rect 880 22912 311728 23192
rect 800 22104 311728 22912
rect 880 21824 311728 22104
rect 800 21152 311728 21824
rect 880 20872 311728 21152
rect 800 20064 311728 20872
rect 880 19784 311728 20064
rect 800 18976 311728 19784
rect 880 18696 311728 18976
rect 800 17888 311728 18696
rect 880 17608 311728 17888
rect 800 16800 311728 17608
rect 880 16520 311728 16800
rect 800 15712 311728 16520
rect 880 15432 311728 15712
rect 800 14624 311728 15432
rect 880 14344 311728 14624
rect 800 13536 311728 14344
rect 880 13256 311728 13536
rect 800 12448 311728 13256
rect 880 12168 311728 12448
rect 800 11360 311728 12168
rect 880 11080 311728 11360
rect 800 10272 311728 11080
rect 880 9992 311728 10272
rect 800 9184 311728 9992
rect 880 8904 311728 9184
rect 800 8096 311728 8904
rect 880 7816 311728 8096
rect 800 7008 311728 7816
rect 880 6728 311728 7008
rect 800 5920 311728 6728
rect 880 5640 311728 5920
rect 800 4832 311728 5640
rect 880 4552 311728 4832
rect 800 3744 311728 4552
rect 880 3464 311728 3744
rect 800 2656 311728 3464
rect 880 2376 311728 2656
rect 800 1568 311728 2376
rect 880 1288 311728 1568
rect 800 616 311728 1288
rect 880 443 311728 616
<< metal4 >>
rect 4208 2128 4528 317744
rect 19568 2128 19888 317744
rect 34928 2128 35248 317744
rect 50288 2128 50608 317744
rect 65648 2128 65968 317744
rect 81008 2128 81328 317744
rect 96368 2128 96688 317744
rect 111728 2128 112048 317744
rect 127088 2128 127408 317744
rect 142448 2128 142768 317744
rect 157808 2128 158128 317744
rect 173168 2128 173488 317744
rect 188528 2128 188848 317744
rect 203888 2128 204208 317744
rect 219248 2128 219568 317744
rect 234608 2128 234928 317744
rect 249968 2128 250288 317744
rect 265328 2128 265648 317744
rect 280688 2128 281008 317744
rect 296048 2128 296368 317744
rect 311408 2128 311728 317744
<< obsm4 >>
rect 979 2483 4128 317525
rect 4608 2483 19488 317525
rect 19968 2483 34848 317525
rect 35328 2483 50208 317525
rect 50688 2483 65568 317525
rect 66048 2483 80928 317525
rect 81408 2483 96288 317525
rect 96768 2483 111648 317525
rect 112128 2483 127008 317525
rect 127488 2483 142368 317525
rect 142848 2483 157728 317525
rect 158208 2483 168853 317525
<< labels >>
rlabel metal3 s 0 143080 800 143200 6 bb_addr0[0]
port 1 nsew signal output
rlabel metal3 s 0 201424 800 201544 6 bb_addr0[10]
port 2 nsew signal output
rlabel metal3 s 0 206864 800 206984 6 bb_addr0[11]
port 3 nsew signal output
rlabel metal3 s 0 212304 800 212424 6 bb_addr0[12]
port 4 nsew signal output
rlabel metal3 s 0 217608 800 217728 6 bb_addr0[13]
port 5 nsew signal output
rlabel metal3 s 0 223048 800 223168 6 bb_addr0[14]
port 6 nsew signal output
rlabel metal3 s 0 228488 800 228608 6 bb_addr0[15]
port 7 nsew signal output
rlabel metal3 s 0 233928 800 234048 6 bb_addr0[16]
port 8 nsew signal output
rlabel metal3 s 0 239232 800 239352 6 bb_addr0[17]
port 9 nsew signal output
rlabel metal3 s 0 244672 800 244792 6 bb_addr0[18]
port 10 nsew signal output
rlabel metal3 s 0 250112 800 250232 6 bb_addr0[19]
port 11 nsew signal output
rlabel metal3 s 0 149608 800 149728 6 bb_addr0[1]
port 12 nsew signal output
rlabel metal3 s 0 255552 800 255672 6 bb_addr0[20]
port 13 nsew signal output
rlabel metal3 s 0 260856 800 260976 6 bb_addr0[21]
port 14 nsew signal output
rlabel metal3 s 0 266296 800 266416 6 bb_addr0[22]
port 15 nsew signal output
rlabel metal3 s 0 271736 800 271856 6 bb_addr0[23]
port 16 nsew signal output
rlabel metal3 s 0 277176 800 277296 6 bb_addr0[24]
port 17 nsew signal output
rlabel metal3 s 0 282480 800 282600 6 bb_addr0[25]
port 18 nsew signal output
rlabel metal3 s 0 287920 800 288040 6 bb_addr0[26]
port 19 nsew signal output
rlabel metal3 s 0 293360 800 293480 6 bb_addr0[27]
port 20 nsew signal output
rlabel metal3 s 0 298800 800 298920 6 bb_addr0[28]
port 21 nsew signal output
rlabel metal3 s 0 304104 800 304224 6 bb_addr0[29]
port 22 nsew signal output
rlabel metal3 s 0 156000 800 156120 6 bb_addr0[2]
port 23 nsew signal output
rlabel metal3 s 0 309544 800 309664 6 bb_addr0[30]
port 24 nsew signal output
rlabel metal3 s 0 314984 800 315104 6 bb_addr0[31]
port 25 nsew signal output
rlabel metal3 s 0 162528 800 162648 6 bb_addr0[3]
port 26 nsew signal output
rlabel metal3 s 0 169056 800 169176 6 bb_addr0[4]
port 27 nsew signal output
rlabel metal3 s 0 174360 800 174480 6 bb_addr0[5]
port 28 nsew signal output
rlabel metal3 s 0 179800 800 179920 6 bb_addr0[6]
port 29 nsew signal output
rlabel metal3 s 0 185240 800 185360 6 bb_addr0[7]
port 30 nsew signal output
rlabel metal3 s 0 190680 800 190800 6 bb_addr0[8]
port 31 nsew signal output
rlabel metal3 s 0 195984 800 196104 6 bb_addr0[9]
port 32 nsew signal output
rlabel metal3 s 0 144168 800 144288 6 bb_addr1[0]
port 33 nsew signal output
rlabel metal3 s 0 202512 800 202632 6 bb_addr1[10]
port 34 nsew signal output
rlabel metal3 s 0 207952 800 208072 6 bb_addr1[11]
port 35 nsew signal output
rlabel metal3 s 0 213392 800 213512 6 bb_addr1[12]
port 36 nsew signal output
rlabel metal3 s 0 218696 800 218816 6 bb_addr1[13]
port 37 nsew signal output
rlabel metal3 s 0 224136 800 224256 6 bb_addr1[14]
port 38 nsew signal output
rlabel metal3 s 0 229576 800 229696 6 bb_addr1[15]
port 39 nsew signal output
rlabel metal3 s 0 235016 800 235136 6 bb_addr1[16]
port 40 nsew signal output
rlabel metal3 s 0 240320 800 240440 6 bb_addr1[17]
port 41 nsew signal output
rlabel metal3 s 0 245760 800 245880 6 bb_addr1[18]
port 42 nsew signal output
rlabel metal3 s 0 251200 800 251320 6 bb_addr1[19]
port 43 nsew signal output
rlabel metal3 s 0 150560 800 150680 6 bb_addr1[1]
port 44 nsew signal output
rlabel metal3 s 0 256504 800 256624 6 bb_addr1[20]
port 45 nsew signal output
rlabel metal3 s 0 261944 800 262064 6 bb_addr1[21]
port 46 nsew signal output
rlabel metal3 s 0 267384 800 267504 6 bb_addr1[22]
port 47 nsew signal output
rlabel metal3 s 0 272824 800 272944 6 bb_addr1[23]
port 48 nsew signal output
rlabel metal3 s 0 278128 800 278248 6 bb_addr1[24]
port 49 nsew signal output
rlabel metal3 s 0 283568 800 283688 6 bb_addr1[25]
port 50 nsew signal output
rlabel metal3 s 0 289008 800 289128 6 bb_addr1[26]
port 51 nsew signal output
rlabel metal3 s 0 294448 800 294568 6 bb_addr1[27]
port 52 nsew signal output
rlabel metal3 s 0 299752 800 299872 6 bb_addr1[28]
port 53 nsew signal output
rlabel metal3 s 0 305192 800 305312 6 bb_addr1[29]
port 54 nsew signal output
rlabel metal3 s 0 157088 800 157208 6 bb_addr1[2]
port 55 nsew signal output
rlabel metal3 s 0 310632 800 310752 6 bb_addr1[30]
port 56 nsew signal output
rlabel metal3 s 0 316072 800 316192 6 bb_addr1[31]
port 57 nsew signal output
rlabel metal3 s 0 163616 800 163736 6 bb_addr1[3]
port 58 nsew signal output
rlabel metal3 s 0 170144 800 170264 6 bb_addr1[4]
port 59 nsew signal output
rlabel metal3 s 0 175448 800 175568 6 bb_addr1[5]
port 60 nsew signal output
rlabel metal3 s 0 180888 800 181008 6 bb_addr1[6]
port 61 nsew signal output
rlabel metal3 s 0 186328 800 186448 6 bb_addr1[7]
port 62 nsew signal output
rlabel metal3 s 0 191768 800 191888 6 bb_addr1[8]
port 63 nsew signal output
rlabel metal3 s 0 197072 800 197192 6 bb_addr1[9]
port 64 nsew signal output
rlabel metal3 s 0 139816 800 139936 6 bb_csb0
port 65 nsew signal output
rlabel metal3 s 0 140904 800 141024 6 bb_csb1
port 66 nsew signal output
rlabel metal3 s 0 145256 800 145376 6 bb_din0[0]
port 67 nsew signal output
rlabel metal3 s 0 203600 800 203720 6 bb_din0[10]
port 68 nsew signal output
rlabel metal3 s 0 209040 800 209160 6 bb_din0[11]
port 69 nsew signal output
rlabel metal3 s 0 214344 800 214464 6 bb_din0[12]
port 70 nsew signal output
rlabel metal3 s 0 219784 800 219904 6 bb_din0[13]
port 71 nsew signal output
rlabel metal3 s 0 225224 800 225344 6 bb_din0[14]
port 72 nsew signal output
rlabel metal3 s 0 230664 800 230784 6 bb_din0[15]
port 73 nsew signal output
rlabel metal3 s 0 235968 800 236088 6 bb_din0[16]
port 74 nsew signal output
rlabel metal3 s 0 241408 800 241528 6 bb_din0[17]
port 75 nsew signal output
rlabel metal3 s 0 246848 800 246968 6 bb_din0[18]
port 76 nsew signal output
rlabel metal3 s 0 252288 800 252408 6 bb_din0[19]
port 77 nsew signal output
rlabel metal3 s 0 151648 800 151768 6 bb_din0[1]
port 78 nsew signal output
rlabel metal3 s 0 257592 800 257712 6 bb_din0[20]
port 79 nsew signal output
rlabel metal3 s 0 263032 800 263152 6 bb_din0[21]
port 80 nsew signal output
rlabel metal3 s 0 268472 800 268592 6 bb_din0[22]
port 81 nsew signal output
rlabel metal3 s 0 273912 800 274032 6 bb_din0[23]
port 82 nsew signal output
rlabel metal3 s 0 279216 800 279336 6 bb_din0[24]
port 83 nsew signal output
rlabel metal3 s 0 284656 800 284776 6 bb_din0[25]
port 84 nsew signal output
rlabel metal3 s 0 290096 800 290216 6 bb_din0[26]
port 85 nsew signal output
rlabel metal3 s 0 295536 800 295656 6 bb_din0[27]
port 86 nsew signal output
rlabel metal3 s 0 300840 800 300960 6 bb_din0[28]
port 87 nsew signal output
rlabel metal3 s 0 306280 800 306400 6 bb_din0[29]
port 88 nsew signal output
rlabel metal3 s 0 158176 800 158296 6 bb_din0[2]
port 89 nsew signal output
rlabel metal3 s 0 311720 800 311840 6 bb_din0[30]
port 90 nsew signal output
rlabel metal3 s 0 317160 800 317280 6 bb_din0[31]
port 91 nsew signal output
rlabel metal3 s 0 164704 800 164824 6 bb_din0[3]
port 92 nsew signal output
rlabel metal3 s 0 171096 800 171216 6 bb_din0[4]
port 93 nsew signal output
rlabel metal3 s 0 176536 800 176656 6 bb_din0[5]
port 94 nsew signal output
rlabel metal3 s 0 181976 800 182096 6 bb_din0[6]
port 95 nsew signal output
rlabel metal3 s 0 187416 800 187536 6 bb_din0[7]
port 96 nsew signal output
rlabel metal3 s 0 192720 800 192840 6 bb_din0[8]
port 97 nsew signal output
rlabel metal3 s 0 198160 800 198280 6 bb_din0[9]
port 98 nsew signal output
rlabel metal3 s 0 146344 800 146464 6 bb_dout0[0]
port 99 nsew signal input
rlabel metal3 s 0 204688 800 204808 6 bb_dout0[10]
port 100 nsew signal input
rlabel metal3 s 0 210128 800 210248 6 bb_dout0[11]
port 101 nsew signal input
rlabel metal3 s 0 215432 800 215552 6 bb_dout0[12]
port 102 nsew signal input
rlabel metal3 s 0 220872 800 220992 6 bb_dout0[13]
port 103 nsew signal input
rlabel metal3 s 0 226312 800 226432 6 bb_dout0[14]
port 104 nsew signal input
rlabel metal3 s 0 231752 800 231872 6 bb_dout0[15]
port 105 nsew signal input
rlabel metal3 s 0 237056 800 237176 6 bb_dout0[16]
port 106 nsew signal input
rlabel metal3 s 0 242496 800 242616 6 bb_dout0[17]
port 107 nsew signal input
rlabel metal3 s 0 247936 800 248056 6 bb_dout0[18]
port 108 nsew signal input
rlabel metal3 s 0 253376 800 253496 6 bb_dout0[19]
port 109 nsew signal input
rlabel metal3 s 0 152736 800 152856 6 bb_dout0[1]
port 110 nsew signal input
rlabel metal3 s 0 258680 800 258800 6 bb_dout0[20]
port 111 nsew signal input
rlabel metal3 s 0 264120 800 264240 6 bb_dout0[21]
port 112 nsew signal input
rlabel metal3 s 0 269560 800 269680 6 bb_dout0[22]
port 113 nsew signal input
rlabel metal3 s 0 275000 800 275120 6 bb_dout0[23]
port 114 nsew signal input
rlabel metal3 s 0 280304 800 280424 6 bb_dout0[24]
port 115 nsew signal input
rlabel metal3 s 0 285744 800 285864 6 bb_dout0[25]
port 116 nsew signal input
rlabel metal3 s 0 291184 800 291304 6 bb_dout0[26]
port 117 nsew signal input
rlabel metal3 s 0 296624 800 296744 6 bb_dout0[27]
port 118 nsew signal input
rlabel metal3 s 0 301928 800 302048 6 bb_dout0[28]
port 119 nsew signal input
rlabel metal3 s 0 307368 800 307488 6 bb_dout0[29]
port 120 nsew signal input
rlabel metal3 s 0 159264 800 159384 6 bb_dout0[2]
port 121 nsew signal input
rlabel metal3 s 0 312808 800 312928 6 bb_dout0[30]
port 122 nsew signal input
rlabel metal3 s 0 318248 800 318368 6 bb_dout0[31]
port 123 nsew signal input
rlabel metal3 s 0 165792 800 165912 6 bb_dout0[3]
port 124 nsew signal input
rlabel metal3 s 0 172184 800 172304 6 bb_dout0[4]
port 125 nsew signal input
rlabel metal3 s 0 177624 800 177744 6 bb_dout0[5]
port 126 nsew signal input
rlabel metal3 s 0 183064 800 183184 6 bb_dout0[6]
port 127 nsew signal input
rlabel metal3 s 0 188504 800 188624 6 bb_dout0[7]
port 128 nsew signal input
rlabel metal3 s 0 193808 800 193928 6 bb_dout0[8]
port 129 nsew signal input
rlabel metal3 s 0 199248 800 199368 6 bb_dout0[9]
port 130 nsew signal input
rlabel metal3 s 0 147432 800 147552 6 bb_dout1[0]
port 131 nsew signal input
rlabel metal3 s 0 205776 800 205896 6 bb_dout1[10]
port 132 nsew signal input
rlabel metal3 s 0 211216 800 211336 6 bb_dout1[11]
port 133 nsew signal input
rlabel metal3 s 0 216520 800 216640 6 bb_dout1[12]
port 134 nsew signal input
rlabel metal3 s 0 221960 800 222080 6 bb_dout1[13]
port 135 nsew signal input
rlabel metal3 s 0 227400 800 227520 6 bb_dout1[14]
port 136 nsew signal input
rlabel metal3 s 0 232840 800 232960 6 bb_dout1[15]
port 137 nsew signal input
rlabel metal3 s 0 238144 800 238264 6 bb_dout1[16]
port 138 nsew signal input
rlabel metal3 s 0 243584 800 243704 6 bb_dout1[17]
port 139 nsew signal input
rlabel metal3 s 0 249024 800 249144 6 bb_dout1[18]
port 140 nsew signal input
rlabel metal3 s 0 254464 800 254584 6 bb_dout1[19]
port 141 nsew signal input
rlabel metal3 s 0 153824 800 153944 6 bb_dout1[1]
port 142 nsew signal input
rlabel metal3 s 0 259768 800 259888 6 bb_dout1[20]
port 143 nsew signal input
rlabel metal3 s 0 265208 800 265328 6 bb_dout1[21]
port 144 nsew signal input
rlabel metal3 s 0 270648 800 270768 6 bb_dout1[22]
port 145 nsew signal input
rlabel metal3 s 0 276088 800 276208 6 bb_dout1[23]
port 146 nsew signal input
rlabel metal3 s 0 281392 800 281512 6 bb_dout1[24]
port 147 nsew signal input
rlabel metal3 s 0 286832 800 286952 6 bb_dout1[25]
port 148 nsew signal input
rlabel metal3 s 0 292272 800 292392 6 bb_dout1[26]
port 149 nsew signal input
rlabel metal3 s 0 297712 800 297832 6 bb_dout1[27]
port 150 nsew signal input
rlabel metal3 s 0 303016 800 303136 6 bb_dout1[28]
port 151 nsew signal input
rlabel metal3 s 0 308456 800 308576 6 bb_dout1[29]
port 152 nsew signal input
rlabel metal3 s 0 160352 800 160472 6 bb_dout1[2]
port 153 nsew signal input
rlabel metal3 s 0 313896 800 314016 6 bb_dout1[30]
port 154 nsew signal input
rlabel metal3 s 0 319336 800 319456 6 bb_dout1[31]
port 155 nsew signal input
rlabel metal3 s 0 166880 800 167000 6 bb_dout1[3]
port 156 nsew signal input
rlabel metal3 s 0 173272 800 173392 6 bb_dout1[4]
port 157 nsew signal input
rlabel metal3 s 0 178712 800 178832 6 bb_dout1[5]
port 158 nsew signal input
rlabel metal3 s 0 184152 800 184272 6 bb_dout1[6]
port 159 nsew signal input
rlabel metal3 s 0 189592 800 189712 6 bb_dout1[7]
port 160 nsew signal input
rlabel metal3 s 0 194896 800 195016 6 bb_dout1[8]
port 161 nsew signal input
rlabel metal3 s 0 200336 800 200456 6 bb_dout1[9]
port 162 nsew signal input
rlabel metal3 s 0 141992 800 142112 6 bb_web0
port 163 nsew signal output
rlabel metal3 s 0 148520 800 148640 6 bb_wmask0[0]
port 164 nsew signal output
rlabel metal3 s 0 154912 800 155032 6 bb_wmask0[1]
port 165 nsew signal output
rlabel metal3 s 0 161440 800 161560 6 bb_wmask0[2]
port 166 nsew signal output
rlabel metal3 s 0 167968 800 168088 6 bb_wmask0[3]
port 167 nsew signal output
rlabel metal2 s 2134 0 2190 800 6 clk_g
port 168 nsew signal input
rlabel metal2 s 19154 0 19210 800 6 io_gecerli
port 169 nsew signal output
rlabel metal2 s 23386 0 23442 800 6 io_oeb[0]
port 170 nsew signal output
rlabel metal2 s 108762 0 108818 800 6 io_oeb[10]
port 171 nsew signal output
rlabel metal2 s 117318 0 117374 800 6 io_oeb[11]
port 172 nsew signal output
rlabel metal2 s 125782 0 125838 800 6 io_oeb[12]
port 173 nsew signal output
rlabel metal2 s 134338 0 134394 800 6 io_oeb[13]
port 174 nsew signal output
rlabel metal2 s 142894 0 142950 800 6 io_oeb[14]
port 175 nsew signal output
rlabel metal2 s 151450 0 151506 800 6 io_oeb[15]
port 176 nsew signal output
rlabel metal2 s 159914 0 159970 800 6 io_oeb[16]
port 177 nsew signal output
rlabel metal2 s 168470 0 168526 800 6 io_oeb[17]
port 178 nsew signal output
rlabel metal2 s 177026 0 177082 800 6 io_oeb[18]
port 179 nsew signal output
rlabel metal2 s 185582 0 185638 800 6 io_oeb[19]
port 180 nsew signal output
rlabel metal2 s 31942 0 31998 800 6 io_oeb[1]
port 181 nsew signal output
rlabel metal2 s 194046 0 194102 800 6 io_oeb[20]
port 182 nsew signal output
rlabel metal2 s 202602 0 202658 800 6 io_oeb[21]
port 183 nsew signal output
rlabel metal2 s 211158 0 211214 800 6 io_oeb[22]
port 184 nsew signal output
rlabel metal2 s 219714 0 219770 800 6 io_oeb[23]
port 185 nsew signal output
rlabel metal2 s 228178 0 228234 800 6 io_oeb[24]
port 186 nsew signal output
rlabel metal2 s 236734 0 236790 800 6 io_oeb[25]
port 187 nsew signal output
rlabel metal2 s 245290 0 245346 800 6 io_oeb[26]
port 188 nsew signal output
rlabel metal2 s 253846 0 253902 800 6 io_oeb[27]
port 189 nsew signal output
rlabel metal2 s 262310 0 262366 800 6 io_oeb[28]
port 190 nsew signal output
rlabel metal2 s 270866 0 270922 800 6 io_oeb[29]
port 191 nsew signal output
rlabel metal2 s 40498 0 40554 800 6 io_oeb[2]
port 192 nsew signal output
rlabel metal2 s 279422 0 279478 800 6 io_oeb[30]
port 193 nsew signal output
rlabel metal2 s 287978 0 288034 800 6 io_oeb[31]
port 194 nsew signal output
rlabel metal2 s 296442 0 296498 800 6 io_oeb[32]
port 195 nsew signal output
rlabel metal2 s 300766 0 300822 800 6 io_oeb[33]
port 196 nsew signal output
rlabel metal2 s 304998 0 305054 800 6 io_oeb[34]
port 197 nsew signal output
rlabel metal2 s 309230 0 309286 800 6 io_oeb[35]
port 198 nsew signal output
rlabel metal2 s 313554 0 313610 800 6 io_oeb[36]
port 199 nsew signal output
rlabel metal2 s 317786 0 317842 800 6 io_oeb[37]
port 200 nsew signal output
rlabel metal2 s 49054 0 49110 800 6 io_oeb[3]
port 201 nsew signal output
rlabel metal2 s 57518 0 57574 800 6 io_oeb[4]
port 202 nsew signal output
rlabel metal2 s 66074 0 66130 800 6 io_oeb[5]
port 203 nsew signal output
rlabel metal2 s 74630 0 74686 800 6 io_oeb[6]
port 204 nsew signal output
rlabel metal2 s 83186 0 83242 800 6 io_oeb[7]
port 205 nsew signal output
rlabel metal2 s 91650 0 91706 800 6 io_oeb[8]
port 206 nsew signal output
rlabel metal2 s 100206 0 100262 800 6 io_oeb[9]
port 207 nsew signal output
rlabel metal2 s 27710 0 27766 800 6 io_ps[0]
port 208 nsew signal output
rlabel metal2 s 112994 0 113050 800 6 io_ps[10]
port 209 nsew signal output
rlabel metal2 s 121550 0 121606 800 6 io_ps[11]
port 210 nsew signal output
rlabel metal2 s 130106 0 130162 800 6 io_ps[12]
port 211 nsew signal output
rlabel metal2 s 138570 0 138626 800 6 io_ps[13]
port 212 nsew signal output
rlabel metal2 s 147126 0 147182 800 6 io_ps[14]
port 213 nsew signal output
rlabel metal2 s 155682 0 155738 800 6 io_ps[15]
port 214 nsew signal output
rlabel metal2 s 164238 0 164294 800 6 io_ps[16]
port 215 nsew signal output
rlabel metal2 s 172702 0 172758 800 6 io_ps[17]
port 216 nsew signal output
rlabel metal2 s 181258 0 181314 800 6 io_ps[18]
port 217 nsew signal output
rlabel metal2 s 189814 0 189870 800 6 io_ps[19]
port 218 nsew signal output
rlabel metal2 s 36174 0 36230 800 6 io_ps[1]
port 219 nsew signal output
rlabel metal2 s 198370 0 198426 800 6 io_ps[20]
port 220 nsew signal output
rlabel metal2 s 206834 0 206890 800 6 io_ps[21]
port 221 nsew signal output
rlabel metal2 s 215390 0 215446 800 6 io_ps[22]
port 222 nsew signal output
rlabel metal2 s 223946 0 224002 800 6 io_ps[23]
port 223 nsew signal output
rlabel metal2 s 232502 0 232558 800 6 io_ps[24]
port 224 nsew signal output
rlabel metal2 s 240966 0 241022 800 6 io_ps[25]
port 225 nsew signal output
rlabel metal2 s 249522 0 249578 800 6 io_ps[26]
port 226 nsew signal output
rlabel metal2 s 258078 0 258134 800 6 io_ps[27]
port 227 nsew signal output
rlabel metal2 s 266634 0 266690 800 6 io_ps[28]
port 228 nsew signal output
rlabel metal2 s 275098 0 275154 800 6 io_ps[29]
port 229 nsew signal output
rlabel metal2 s 44730 0 44786 800 6 io_ps[2]
port 230 nsew signal output
rlabel metal2 s 283654 0 283710 800 6 io_ps[30]
port 231 nsew signal output
rlabel metal2 s 292210 0 292266 800 6 io_ps[31]
port 232 nsew signal output
rlabel metal2 s 53286 0 53342 800 6 io_ps[3]
port 233 nsew signal output
rlabel metal2 s 61842 0 61898 800 6 io_ps[4]
port 234 nsew signal output
rlabel metal2 s 70306 0 70362 800 6 io_ps[5]
port 235 nsew signal output
rlabel metal2 s 78862 0 78918 800 6 io_ps[6]
port 236 nsew signal output
rlabel metal2 s 87418 0 87474 800 6 io_ps[7]
port 237 nsew signal output
rlabel metal2 s 95974 0 96030 800 6 io_ps[8]
port 238 nsew signal output
rlabel metal2 s 104438 0 104494 800 6 io_ps[9]
port 239 nsew signal output
rlabel metal2 s 6366 0 6422 800 6 rst_g
port 240 nsew signal input
rlabel metal2 s 14922 0 14978 800 6 rx
port 241 nsew signal input
rlabel metal2 s 10598 0 10654 800 6 tx
port 242 nsew signal output
rlabel metal3 s 0 3544 800 3664 6 vb_addr0[0]
port 243 nsew signal output
rlabel metal3 s 0 62024 800 62144 6 vb_addr0[10]
port 244 nsew signal output
rlabel metal3 s 0 67328 800 67448 6 vb_addr0[11]
port 245 nsew signal output
rlabel metal3 s 0 72768 800 72888 6 vb_addr0[12]
port 246 nsew signal output
rlabel metal3 s 0 10072 800 10192 6 vb_addr0[1]
port 247 nsew signal output
rlabel metal3 s 0 16600 800 16720 6 vb_addr0[2]
port 248 nsew signal output
rlabel metal3 s 0 22992 800 23112 6 vb_addr0[3]
port 249 nsew signal output
rlabel metal3 s 0 29520 800 29640 6 vb_addr0[4]
port 250 nsew signal output
rlabel metal3 s 0 34960 800 35080 6 vb_addr0[5]
port 251 nsew signal output
rlabel metal3 s 0 40400 800 40520 6 vb_addr0[6]
port 252 nsew signal output
rlabel metal3 s 0 45704 800 45824 6 vb_addr0[7]
port 253 nsew signal output
rlabel metal3 s 0 51144 800 51264 6 vb_addr0[8]
port 254 nsew signal output
rlabel metal3 s 0 56584 800 56704 6 vb_addr0[9]
port 255 nsew signal output
rlabel metal3 s 0 4632 800 4752 6 vb_addr1[0]
port 256 nsew signal output
rlabel metal3 s 0 63112 800 63232 6 vb_addr1[10]
port 257 nsew signal output
rlabel metal3 s 0 68416 800 68536 6 vb_addr1[11]
port 258 nsew signal output
rlabel metal3 s 0 73856 800 73976 6 vb_addr1[12]
port 259 nsew signal output
rlabel metal3 s 0 11160 800 11280 6 vb_addr1[1]
port 260 nsew signal output
rlabel metal3 s 0 17688 800 17808 6 vb_addr1[2]
port 261 nsew signal output
rlabel metal3 s 0 24080 800 24200 6 vb_addr1[3]
port 262 nsew signal output
rlabel metal3 s 0 30608 800 30728 6 vb_addr1[4]
port 263 nsew signal output
rlabel metal3 s 0 36048 800 36168 6 vb_addr1[5]
port 264 nsew signal output
rlabel metal3 s 0 41488 800 41608 6 vb_addr1[6]
port 265 nsew signal output
rlabel metal3 s 0 46792 800 46912 6 vb_addr1[7]
port 266 nsew signal output
rlabel metal3 s 0 52232 800 52352 6 vb_addr1[8]
port 267 nsew signal output
rlabel metal3 s 0 57672 800 57792 6 vb_addr1[9]
port 268 nsew signal output
rlabel metal3 s 0 416 800 536 6 vb_csb0
port 269 nsew signal output
rlabel metal3 s 0 1368 800 1488 6 vb_csb1
port 270 nsew signal output
rlabel metal3 s 0 5720 800 5840 6 vb_din0[0]
port 271 nsew signal output
rlabel metal3 s 0 64200 800 64320 6 vb_din0[10]
port 272 nsew signal output
rlabel metal3 s 0 69504 800 69624 6 vb_din0[11]
port 273 nsew signal output
rlabel metal3 s 0 74944 800 75064 6 vb_din0[12]
port 274 nsew signal output
rlabel metal3 s 0 78208 800 78328 6 vb_din0[13]
port 275 nsew signal output
rlabel metal3 s 0 81472 800 81592 6 vb_din0[14]
port 276 nsew signal output
rlabel metal3 s 0 84736 800 84856 6 vb_din0[15]
port 277 nsew signal output
rlabel metal3 s 0 87864 800 87984 6 vb_din0[16]
port 278 nsew signal output
rlabel metal3 s 0 91128 800 91248 6 vb_din0[17]
port 279 nsew signal output
rlabel metal3 s 0 94392 800 94512 6 vb_din0[18]
port 280 nsew signal output
rlabel metal3 s 0 97656 800 97776 6 vb_din0[19]
port 281 nsew signal output
rlabel metal3 s 0 12248 800 12368 6 vb_din0[1]
port 282 nsew signal output
rlabel metal3 s 0 100920 800 101040 6 vb_din0[20]
port 283 nsew signal output
rlabel metal3 s 0 104184 800 104304 6 vb_din0[21]
port 284 nsew signal output
rlabel metal3 s 0 107312 800 107432 6 vb_din0[22]
port 285 nsew signal output
rlabel metal3 s 0 110576 800 110696 6 vb_din0[23]
port 286 nsew signal output
rlabel metal3 s 0 113840 800 113960 6 vb_din0[24]
port 287 nsew signal output
rlabel metal3 s 0 117104 800 117224 6 vb_din0[25]
port 288 nsew signal output
rlabel metal3 s 0 120368 800 120488 6 vb_din0[26]
port 289 nsew signal output
rlabel metal3 s 0 123632 800 123752 6 vb_din0[27]
port 290 nsew signal output
rlabel metal3 s 0 126896 800 127016 6 vb_din0[28]
port 291 nsew signal output
rlabel metal3 s 0 130024 800 130144 6 vb_din0[29]
port 292 nsew signal output
rlabel metal3 s 0 18776 800 18896 6 vb_din0[2]
port 293 nsew signal output
rlabel metal3 s 0 133288 800 133408 6 vb_din0[30]
port 294 nsew signal output
rlabel metal3 s 0 136552 800 136672 6 vb_din0[31]
port 295 nsew signal output
rlabel metal3 s 0 25168 800 25288 6 vb_din0[3]
port 296 nsew signal output
rlabel metal3 s 0 31696 800 31816 6 vb_din0[4]
port 297 nsew signal output
rlabel metal3 s 0 37136 800 37256 6 vb_din0[5]
port 298 nsew signal output
rlabel metal3 s 0 42576 800 42696 6 vb_din0[6]
port 299 nsew signal output
rlabel metal3 s 0 47880 800 48000 6 vb_din0[7]
port 300 nsew signal output
rlabel metal3 s 0 53320 800 53440 6 vb_din0[8]
port 301 nsew signal output
rlabel metal3 s 0 58760 800 58880 6 vb_din0[9]
port 302 nsew signal output
rlabel metal3 s 0 6808 800 6928 6 vb_dout0[0]
port 303 nsew signal input
rlabel metal3 s 0 65152 800 65272 6 vb_dout0[10]
port 304 nsew signal input
rlabel metal3 s 0 70592 800 70712 6 vb_dout0[11]
port 305 nsew signal input
rlabel metal3 s 0 76032 800 76152 6 vb_dout0[12]
port 306 nsew signal input
rlabel metal3 s 0 79296 800 79416 6 vb_dout0[13]
port 307 nsew signal input
rlabel metal3 s 0 82560 800 82680 6 vb_dout0[14]
port 308 nsew signal input
rlabel metal3 s 0 85688 800 85808 6 vb_dout0[15]
port 309 nsew signal input
rlabel metal3 s 0 88952 800 89072 6 vb_dout0[16]
port 310 nsew signal input
rlabel metal3 s 0 92216 800 92336 6 vb_dout0[17]
port 311 nsew signal input
rlabel metal3 s 0 95480 800 95600 6 vb_dout0[18]
port 312 nsew signal input
rlabel metal3 s 0 98744 800 98864 6 vb_dout0[19]
port 313 nsew signal input
rlabel metal3 s 0 13336 800 13456 6 vb_dout0[1]
port 314 nsew signal input
rlabel metal3 s 0 102008 800 102128 6 vb_dout0[20]
port 315 nsew signal input
rlabel metal3 s 0 105272 800 105392 6 vb_dout0[21]
port 316 nsew signal input
rlabel metal3 s 0 108400 800 108520 6 vb_dout0[22]
port 317 nsew signal input
rlabel metal3 s 0 111664 800 111784 6 vb_dout0[23]
port 318 nsew signal input
rlabel metal3 s 0 114928 800 115048 6 vb_dout0[24]
port 319 nsew signal input
rlabel metal3 s 0 118192 800 118312 6 vb_dout0[25]
port 320 nsew signal input
rlabel metal3 s 0 121456 800 121576 6 vb_dout0[26]
port 321 nsew signal input
rlabel metal3 s 0 124720 800 124840 6 vb_dout0[27]
port 322 nsew signal input
rlabel metal3 s 0 127984 800 128104 6 vb_dout0[28]
port 323 nsew signal input
rlabel metal3 s 0 131112 800 131232 6 vb_dout0[29]
port 324 nsew signal input
rlabel metal3 s 0 19864 800 19984 6 vb_dout0[2]
port 325 nsew signal input
rlabel metal3 s 0 134376 800 134496 6 vb_dout0[30]
port 326 nsew signal input
rlabel metal3 s 0 137640 800 137760 6 vb_dout0[31]
port 327 nsew signal input
rlabel metal3 s 0 26256 800 26376 6 vb_dout0[3]
port 328 nsew signal input
rlabel metal3 s 0 32784 800 32904 6 vb_dout0[4]
port 329 nsew signal input
rlabel metal3 s 0 38224 800 38344 6 vb_dout0[5]
port 330 nsew signal input
rlabel metal3 s 0 43528 800 43648 6 vb_dout0[6]
port 331 nsew signal input
rlabel metal3 s 0 48968 800 49088 6 vb_dout0[7]
port 332 nsew signal input
rlabel metal3 s 0 54408 800 54528 6 vb_dout0[8]
port 333 nsew signal input
rlabel metal3 s 0 59848 800 59968 6 vb_dout0[9]
port 334 nsew signal input
rlabel metal3 s 0 7896 800 8016 6 vb_dout1[0]
port 335 nsew signal input
rlabel metal3 s 0 66240 800 66360 6 vb_dout1[10]
port 336 nsew signal input
rlabel metal3 s 0 71680 800 71800 6 vb_dout1[11]
port 337 nsew signal input
rlabel metal3 s 0 77120 800 77240 6 vb_dout1[12]
port 338 nsew signal input
rlabel metal3 s 0 80384 800 80504 6 vb_dout1[13]
port 339 nsew signal input
rlabel metal3 s 0 83648 800 83768 6 vb_dout1[14]
port 340 nsew signal input
rlabel metal3 s 0 86776 800 86896 6 vb_dout1[15]
port 341 nsew signal input
rlabel metal3 s 0 90040 800 90160 6 vb_dout1[16]
port 342 nsew signal input
rlabel metal3 s 0 93304 800 93424 6 vb_dout1[17]
port 343 nsew signal input
rlabel metal3 s 0 96568 800 96688 6 vb_dout1[18]
port 344 nsew signal input
rlabel metal3 s 0 99832 800 99952 6 vb_dout1[19]
port 345 nsew signal input
rlabel metal3 s 0 14424 800 14544 6 vb_dout1[1]
port 346 nsew signal input
rlabel metal3 s 0 103096 800 103216 6 vb_dout1[20]
port 347 nsew signal input
rlabel metal3 s 0 106360 800 106480 6 vb_dout1[21]
port 348 nsew signal input
rlabel metal3 s 0 109488 800 109608 6 vb_dout1[22]
port 349 nsew signal input
rlabel metal3 s 0 112752 800 112872 6 vb_dout1[23]
port 350 nsew signal input
rlabel metal3 s 0 116016 800 116136 6 vb_dout1[24]
port 351 nsew signal input
rlabel metal3 s 0 119280 800 119400 6 vb_dout1[25]
port 352 nsew signal input
rlabel metal3 s 0 122544 800 122664 6 vb_dout1[26]
port 353 nsew signal input
rlabel metal3 s 0 125808 800 125928 6 vb_dout1[27]
port 354 nsew signal input
rlabel metal3 s 0 128936 800 129056 6 vb_dout1[28]
port 355 nsew signal input
rlabel metal3 s 0 132200 800 132320 6 vb_dout1[29]
port 356 nsew signal input
rlabel metal3 s 0 20952 800 21072 6 vb_dout1[2]
port 357 nsew signal input
rlabel metal3 s 0 135464 800 135584 6 vb_dout1[30]
port 358 nsew signal input
rlabel metal3 s 0 138728 800 138848 6 vb_dout1[31]
port 359 nsew signal input
rlabel metal3 s 0 27344 800 27464 6 vb_dout1[3]
port 360 nsew signal input
rlabel metal3 s 0 33872 800 33992 6 vb_dout1[4]
port 361 nsew signal input
rlabel metal3 s 0 39312 800 39432 6 vb_dout1[5]
port 362 nsew signal input
rlabel metal3 s 0 44616 800 44736 6 vb_dout1[6]
port 363 nsew signal input
rlabel metal3 s 0 50056 800 50176 6 vb_dout1[7]
port 364 nsew signal input
rlabel metal3 s 0 55496 800 55616 6 vb_dout1[8]
port 365 nsew signal input
rlabel metal3 s 0 60936 800 61056 6 vb_dout1[9]
port 366 nsew signal input
rlabel metal3 s 0 2456 800 2576 6 vb_web0
port 367 nsew signal output
rlabel metal3 s 0 8984 800 9104 6 vb_wmask0[0]
port 368 nsew signal output
rlabel metal3 s 0 15512 800 15632 6 vb_wmask0[1]
port 369 nsew signal output
rlabel metal3 s 0 21904 800 22024 6 vb_wmask0[2]
port 370 nsew signal output
rlabel metal3 s 0 28432 800 28552 6 vb_wmask0[3]
port 371 nsew signal output
rlabel metal4 s 4208 2128 4528 317744 6 vccd1
port 372 nsew power input
rlabel metal4 s 34928 2128 35248 317744 6 vccd1
port 372 nsew power input
rlabel metal4 s 65648 2128 65968 317744 6 vccd1
port 372 nsew power input
rlabel metal4 s 96368 2128 96688 317744 6 vccd1
port 372 nsew power input
rlabel metal4 s 127088 2128 127408 317744 6 vccd1
port 372 nsew power input
rlabel metal4 s 157808 2128 158128 317744 6 vccd1
port 372 nsew power input
rlabel metal4 s 188528 2128 188848 317744 6 vccd1
port 372 nsew power input
rlabel metal4 s 219248 2128 219568 317744 6 vccd1
port 372 nsew power input
rlabel metal4 s 249968 2128 250288 317744 6 vccd1
port 372 nsew power input
rlabel metal4 s 280688 2128 281008 317744 6 vccd1
port 372 nsew power input
rlabel metal4 s 311408 2128 311728 317744 6 vccd1
port 372 nsew power input
rlabel metal4 s 19568 2128 19888 317744 6 vssd1
port 373 nsew ground input
rlabel metal4 s 50288 2128 50608 317744 6 vssd1
port 373 nsew ground input
rlabel metal4 s 81008 2128 81328 317744 6 vssd1
port 373 nsew ground input
rlabel metal4 s 111728 2128 112048 317744 6 vssd1
port 373 nsew ground input
rlabel metal4 s 142448 2128 142768 317744 6 vssd1
port 373 nsew ground input
rlabel metal4 s 173168 2128 173488 317744 6 vssd1
port 373 nsew ground input
rlabel metal4 s 203888 2128 204208 317744 6 vssd1
port 373 nsew ground input
rlabel metal4 s 234608 2128 234928 317744 6 vssd1
port 373 nsew ground input
rlabel metal4 s 265328 2128 265648 317744 6 vssd1
port 373 nsew ground input
rlabel metal4 s 296048 2128 296368 317744 6 vssd1
port 373 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 320000 320000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 79676308
string GDS_FILE /home/kasirga/c0_hayyan/GL_GECTI/caravel_user_project/openlane/c0_system/runs/c0_system/results/finishing/c0_system.magic.gds
string GDS_START 1683532
<< end >>

